library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.TIPOS.all;

entity paddle1 is
	port(
		--Essential
		clk, reset:				 in std_logic;
		pixel_x, pixel_y:		 in std_logic_vector(9 downto 0);
		stop_game:				 in std_logic;
		
		--Reset Position with Score
		goal_tick:				 in std_logic_vector(1 downto 0);
		
		--Joystick
		refresh_tick_pad:		 in std_logic;
		pad1_Ry_EN:				 in std_logic;
		pad1_Ry:					 in std_logic;
		pad1_Rx_EN:				 in std_logic;
		pad1_Rx:					 in std_logic;
				
		--Pad Position
		pad_X:					out std_logic_vector(9 downto 0);
		pad_Y:					out std_logic_vector(9 downto 0);
		
		--Pad Video Information
		obj_on:				out std_logic;
		obj_RGB:				out TYPE_COR
	);
	
end paddle1;

architecture arch of paddle1 is
	signal forced_rst: std_logic := '0';
	
	--Definicoes basicas da img
	constant LINHAS:  integer := 61;
   constant COLUNAS: integer := 61;
	constant N_CORES:	integer := 30;
	--Dimensoes da Imagem na tela
	signal obj_Ymin: integer := (480-LINHAS)/2;
	signal obj_Xmin: integer := 50;
	signal obj_Ymax: integer := obj_Ymin + LINHAS;
	signal obj_Xmax: integer := obj_Xmin + COLUNAS;
	
	signal obj_Ymin_next: integer := obj_Ymin;
	signal obj_Xmin_next: integer := obj_Xmin;
	
	constant frontier_Xmax: integer := 640 - 25 - COLUNAS;
	constant frontier_Xmin: integer := 318;
	constant frontier_Ymin: integer := 26  + 15;
	constant frontier_Ymax: integer := 454 - 13 - LINHAS;
	--Definindo a img
	type linha_bitmap is array(0 to COLUNAS -1) of integer range 0 to N_CORES;
	type   obj_bitmap is array(0 to LINHAS  -1) of linha_bitmap;
	
   constant obj_matriz: obj_bitmap :=
	(
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3, 3, 2, 2, 1, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 6, 7, 3, 8, 8, 8, 8, 8, 8, 8, 9, 8, 8, 8, 8, 8, 8, 8, 7, 6, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 11, 12, 13, 8, 8, 9, 14, 14, 15, 15, 15, 15, 15, 15, 16, 17, 14, 14, 9, 9, 8, 13, 12, 11, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 11, 12, 13, 8, 18, 15, 15, 16, 16, 19, 19, 19, 16, 16, 16, 16, 16, 16, 16, 20, 20, 20, 17, 18, 8, 13, 12, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 6, 12, 13, 8, 17, 20, 16, 15, 15, 16, 20, 19, 19, 20, 20, 20, 19, 20, 20, 20, 21, 21, 21, 21, 21, 19, 17, 14, 8, 13, 12, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 11, 13, 8, 9, 17, 20, 21, 19, 19, 16, 16, 20, 20, 20, 20, 20, 21, 21, 20, 20, 20, 20, 20, 20, 20, 20, 19, 20, 19, 20, 18, 8, 13, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 7, 8, 18, 17, 16, 19, 16, 20, 19, 21, 20, 20, 16, 20, 17, 17, 17, 17, 17, 14, 17, 16, 15, 16, 16, 19, 19, 20, 16, 15, 16, 19, 14, 9, 13, 7, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 12, 8, 9, 21, 20, 16, 16, 15, 15, 16, 20, 17, 17, 14, 9, 9, 9, 8, 8, 8, 8, 9, 9, 14, 14, 14, 20, 19, 20, 16, 15, 15, 16, 19, 20, 9, 13, 12, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 12, 8, 14, 16, 20, 20, 16, 16, 15, 15, 15, 17, 18, 8, 8, 13, 13, 22, 22, 22, 22, 22, 13, 13, 13, 8, 18, 18, 17, 20, 20, 16, 16, 16, 16, 20, 16, 14, 8, 12, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 10, 12, 8, 17, 20, 19, 16, 16, 20, 19, 20, 14, 18, 8, 13, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 13, 13, 8, 18, 17, 20, 19, 16, 16, 16, 16, 20, 17, 8, 12, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 5, 12, 13, 17, 21, 15, 16, 16, 20, 19, 20, 17, 18, 13, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 13, 18, 17, 20, 16, 16, 15, 16, 16, 16, 14, 13, 12, 5, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 4, 11, 8, 14, 21, 16, 15, 16, 16, 20, 17, 18, 8, 13, 22, 22, 22, 22, 22, 22, 13, 13, 13, 13, 13, 13, 13, 13, 22, 22, 22, 22, 22, 22, 13, 8, 14, 20, 16, 15, 16, 19, 16, 16, 17, 13, 7, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 6, 13, 14, 19, 19, 15, 16, 19, 20, 17, 18, 13, 22, 22, 22, 22, 13, 13, 13, 13, 8, 8, 8, 8, 8, 8, 8, 8, 13, 13, 13, 22, 22, 22, 22, 22, 8, 18, 17, 19, 19, 19, 15, 15, 19, 18, 12, 11, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 10, 12, 8, 15, 16, 16, 16, 16, 20, 17, 18, 13, 22, 22, 22, 22, 13, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 13, 22, 22, 22, 22, 8, 18, 20, 19, 20, 15, 16, 19, 17, 18, 18, 5, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 7, 8, 21, 20, 16, 16, 16, 16, 17, 14, 13, 22, 22, 22, 13, 13, 8, 8, 8, 8, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 8, 8, 8, 13, 13, 22, 22, 22, 8, 14, 20, 21, 20, 19, 20, 20, 17, 9, 11, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 6, 12, 14, 19, 20, 16, 16, 20, 20, 17, 8, 22, 22, 22, 13, 8, 8, 8, 9, 18, 18, 18, 18, 18, 14, 14, 14, 14, 14, 18, 18, 18, 18, 8, 8, 8, 13, 13, 22, 22, 22, 8, 18, 21, 21, 16, 16, 19, 15, 14, 12, 6, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 7, 18, 15, 16, 20, 20, 16, 20, 17, 18, 13, 22, 22, 13, 8, 8, 8, 18, 18, 14, 14, 14, 14, 17, 17, 17, 17, 14, 14, 14, 14, 14, 9, 18, 18, 8, 8, 13, 13, 22, 22, 13, 18, 17, 21, 16, 16, 16, 15, 15, 9, 7, 0, 0, 0, 0, 0),
		(0, 0, 0, 10, 12, 17, 20, 20, 20, 19, 19, 20, 18, 13, 22, 13, 13, 8, 8, 18, 18, 18, 14, 14, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 14, 14, 14, 18, 8, 8, 8, 8, 13, 22, 22, 13, 14, 21, 20, 16, 16, 16, 20, 9, 12, 10, 0, 0, 0, 0),
		(0, 0, 0, 11, 8, 17, 20, 16, 15, 16, 19, 17, 8, 13, 22, 13, 8, 8, 18, 18, 18, 14, 17, 17, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 17, 17, 17, 14, 18, 18, 18, 8, 8, 13, 22, 13, 9, 17, 21, 16, 16, 16, 20, 17, 18, 11, 0, 0, 0, 0),
		(0, 0, 5, 12, 18, 20, 20, 16, 15, 16, 20, 18, 13, 13, 13, 8, 8, 18, 18, 14, 17, 17, 17, 20, 16, 20, 20, 19, 19, 19, 20, 19, 16, 20, 20, 20, 20, 17, 17, 14, 14, 18, 8, 8, 8, 22, 22, 8, 17, 21, 20, 16, 16, 20, 21, 17, 12, 5, 0, 0, 0),
		(0, 0, 6, 8, 17, 15, 20, 16, 16, 19, 17, 18, 13, 13, 13, 8, 18, 18, 14, 17, 17, 20, 20, 16, 16, 16, 19, 19, 19, 20, 16, 16, 16, 16, 20, 20, 20, 20, 20, 17, 17, 18, 18, 18, 8, 13, 13, 13, 18, 21, 21, 16, 16, 16, 20, 17, 8, 6, 0, 0, 0),
		(0, 0, 7, 18, 15, 15, 20, 19, 19, 21, 17, 8, 13, 13, 8, 18, 18, 14, 17, 17, 20, 16, 16, 16, 16, 16, 19, 19, 19, 20, 16, 16, 16, 16, 20, 20, 20, 20, 20, 20, 17, 14, 18, 18, 18, 8, 13, 13, 8, 17, 21, 20, 16, 16, 20, 21, 18, 11, 0, 0, 0),
		(0, 4, 12, 17, 15, 15, 16, 20, 16, 20, 18, 13, 13, 13, 8, 18, 14, 17, 17, 20, 16, 15, 15, 16, 20, 16, 20, 20, 20, 16, 16, 16, 16, 20, 20, 20, 20, 20, 20, 16, 17, 17, 17, 18, 18, 8, 8, 13, 13, 14, 21, 20, 16, 16, 19, 20, 14, 12, 0, 0, 0),
		(0, 10, 18, 15, 16, 15, 16, 16, 20, 21, 18, 13, 13, 8, 18, 14, 14, 17, 20, 20, 16, 16, 16, 16, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 17, 14, 18, 18, 8, 13, 13, 18, 17, 16, 16, 20, 16, 16, 17, 12, 10, 0, 0),
		(0, 6, 9, 15, 16, 16, 15, 16, 21, 21, 8, 13, 13, 8, 18, 14, 14, 17, 20, 20, 16, 16, 16, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 17, 14, 14, 9, 9, 13, 13, 18, 17, 15, 19, 21, 16, 16, 16, 18, 6, 0, 0),
		(0, 11, 18, 16, 16, 19, 16, 16, 21, 17, 8, 13, 8, 8, 18, 14, 17, 20, 20, 20, 16, 16, 16, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 17, 17, 14, 18, 9, 8, 13, 8, 17, 15, 19, 21, 20, 16, 16, 18, 6, 0, 0),
		(0, 7, 14, 16, 16, 19, 19, 16, 19, 17, 8, 13, 8, 18, 14, 14, 17, 20, 20, 20, 16, 16, 16, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 16, 16, 20, 20, 20, 17, 14, 14, 18, 8, 13, 8, 17, 16, 19, 21, 20, 16, 16, 18, 11, 0, 0),
		(0, 7, 14, 16, 15, 19, 19, 16, 20, 17, 8, 13, 18, 18, 14, 14, 17, 20, 20, 20, 16, 16, 16, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 16, 16, 16, 20, 20, 17, 17, 14, 14, 8, 13, 8, 17, 16, 16, 20, 21, 16, 16, 17, 7, 0, 0),
		(0, 12, 17, 15, 15, 19, 20, 16, 20, 17, 8, 8, 18, 17, 14, 17, 17, 20, 20, 20, 20, 16, 16, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 16, 16, 16, 19, 20, 20, 17, 14, 14, 18, 13, 8, 17, 16, 16, 20, 20, 16, 15, 17, 12, 0, 0),
		(0, 12, 17, 15, 15, 21, 20, 16, 19, 14, 8, 8, 18, 17, 17, 17, 17, 20, 20, 20, 20, 16, 16, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 16, 16, 16, 16, 20, 20, 17, 17, 14, 18, 8, 8, 17, 16, 16, 20, 17, 16, 15, 17, 12, 0, 0),
		(0, 12, 17, 15, 19, 21, 20, 20, 19, 17, 8, 8, 18, 17, 14, 17, 20, 20, 20, 19, 20, 16, 16, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 16, 15, 16, 16, 20, 20, 17, 14, 14, 18, 8, 8, 17, 15, 15, 20, 17, 16, 15, 17, 12, 0, 0),
		(0, 12, 17, 15, 19, 19, 20, 20, 19, 17, 8, 8, 18, 17, 17, 17, 17, 21, 19, 20, 16, 16, 19, 19, 20, 20, 20, 20, 20, 20, 20, 16, 16, 16, 16, 20, 20, 20, 20, 16, 16, 19, 20, 20, 17, 14, 17, 18, 8, 8, 17, 16, 16, 20, 21, 19, 15, 14, 12, 0, 0),
		(0, 12, 17, 16, 15, 16, 20, 16, 19, 17, 9, 8, 18, 17, 17, 17, 17, 21, 21, 16, 16, 15, 19, 19, 20, 20, 20, 20, 20, 20, 20, 15, 16, 16, 16, 16, 20, 20, 21, 20, 19, 19, 16, 16, 17, 14, 17, 18, 8, 9, 20, 20, 20, 20, 20, 16, 19, 14, 12, 0, 0),
		(0, 7, 17, 15, 15, 19, 20, 16, 19, 20, 9, 8, 18, 17, 17, 21, 17, 21, 23, 21, 19, 16, 16, 20, 20, 20, 20, 20, 20, 20, 20, 19, 16, 16, 16, 16, 20, 20, 19, 21, 21, 23, 19, 16, 17, 14, 17, 18, 8, 9, 21, 20, 20, 20, 20, 16, 16, 17, 7, 0, 0),
		(0, 7, 17, 16, 15, 19, 20, 16, 19, 20, 9, 8, 18, 17, 17, 20, 17, 21, 24, 23, 21, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 16, 16, 16, 16, 20, 20, 20, 20, 21, 23, 23, 19, 17, 17, 14, 14, 18, 8, 14, 21, 20, 20, 20, 20, 16, 16, 17, 11, 0, 0),
		(0, 11, 14, 19, 16, 20, 20, 16, 19, 21, 14, 9, 9, 14, 17, 17, 17, 23, 25, 24, 23, 21, 20, 20, 20, 20, 20, 20, 20, 20, 20, 16, 16, 16, 20, 20, 20, 20, 21, 23, 24, 25, 23, 17, 17, 17, 14, 8, 8, 17, 19, 20, 19, 20, 20, 19, 19, 17, 6, 0, 0),
		(0, 10, 18, 19, 19, 17, 20, 19, 16, 19, 17, 9, 9, 14, 17, 16, 15, 23, 25, 25, 24, 21, 20, 20, 20, 20, 20, 20, 20, 20, 20, 16, 20, 20, 20, 20, 20, 20, 21, 24, 25, 25, 23, 14, 17, 17, 14, 8, 9, 20, 19, 20, 19, 16, 20, 19, 19, 18, 10, 0, 0),
		(0, 5, 12, 19, 21, 20, 20, 19, 16, 20, 20, 14, 9, 9, 14, 16, 16, 23, 25, 26, 25, 24, 21, 20, 19, 19, 20, 20, 20, 20, 20, 19, 19, 20, 20, 20, 21, 23, 24, 25, 26, 25, 21, 14, 17, 14, 9, 8, 14, 21, 20, 20, 16, 16, 20, 23, 21, 12, 4, 0, 0),
		(0, 0, 12, 20, 23, 21, 20, 19, 16, 20, 21, 17, 9, 9, 14, 15, 15, 21, 25, 1, 26, 25, 23, 19, 19, 21, 21, 20, 20, 20, 20, 20, 19, 20, 20, 20, 23, 24, 25, 26, 1, 25, 17, 17, 17, 14, 9, 8, 17, 21, 20, 16, 16, 16, 19, 23, 21, 7, 0, 0, 0),
		(0, 0, 7, 17, 23, 19, 20, 20, 16, 16, 19, 20, 9, 9, 18, 15, 14, 17, 25, 1, 1, 26, 25, 23, 21, 19, 19, 19, 16, 16, 17, 20, 20, 19, 16, 21, 24, 25, 26, 1, 1, 25, 14, 17, 17, 9, 9, 9, 21, 21, 16, 16, 16, 16, 21, 23, 21, 11, 0, 0, 0),
		(0, 0, 10, 12, 19, 19, 19, 20, 19, 16, 16, 16, 14, 9, 18, 17, 14, 14, 24, 1, 27, 27, 1, 25, 24, 21, 16, 15, 15, 15, 20, 17, 20, 19, 21, 24, 25, 1, 27, 27, 26, 23, 15, 15, 17, 18, 9, 15, 19, 20, 20, 16, 16, 16, 23, 23, 12, 10, 0, 0, 0),
		(0, 0, 0, 12, 19, 19, 19, 21, 20, 16, 16, 19, 20, 9, 8, 14, 20, 14, 17, 25, 27, 28, 27, 1, 26, 25, 23, 19, 16, 17, 21, 21, 21, 23, 25, 26, 1, 27, 28, 27, 25, 17, 15, 15, 9, 8, 14, 16, 16, 19, 20, 20, 16, 19, 23, 21, 12, 0, 0, 0, 0),
		(0, 0, 0, 11, 14, 23, 23, 20, 20, 19, 16, 16, 21, 17, 9, 9, 14, 20, 14, 21, 26, 28, 28, 28, 27, 1, 1, 26, 25, 25, 25, 25, 26, 1, 27, 28, 28, 28, 28, 26, 21, 14, 21, 14, 9, 18, 21, 20, 17, 20, 20, 19, 15, 23, 24, 17, 11, 0, 0, 0, 0),
		(0, 0, 0, 5, 12, 24, 24, 21, 20, 19, 16, 16, 19, 21, 17, 8, 9, 17, 16, 17, 24, 1, 28, 29, 29, 29, 28, 28, 28, 28, 28, 28, 28, 28, 29, 29, 29, 28, 1, 21, 14, 17, 21, 18, 9, 21, 21, 16, 20, 17, 20, 20, 20, 24, 23, 12, 5, 0, 0, 0, 0),
		(0, 0, 0, 0, 11, 17, 25, 24, 20, 20, 16, 16, 19, 21, 20, 18, 18, 9, 14, 16, 14, 24, 1, 28, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 28, 1, 24, 15, 14, 17, 18, 18, 17, 21, 20, 16, 20, 20, 20, 17, 24, 25, 18, 11, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 5, 12, 25, 25, 23, 20, 16, 16, 16, 20, 20, 21, 17, 9, 9, 17, 17, 14, 24, 1, 28, 29, 29, 29, 29, 29, 29, 29, 29, 29, 28, 27, 26, 23, 14, 17, 17, 9, 9, 14, 21, 19, 15, 16, 16, 21, 21, 23, 25, 24, 12, 5, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 11, 17, 25, 25, 20, 16, 19, 16, 16, 20, 21, 21, 17, 9, 9, 14, 14, 17, 21, 25, 1, 27, 28, 28, 29, 29, 28, 28, 27, 1, 25, 21, 14, 14, 17, 18, 9, 14, 16, 16, 15, 16, 15, 16, 20, 21, 25, 25, 12, 6, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 4, 12, 24, 26, 23, 15, 15, 21, 21, 19, 20, 19, 21, 17, 9, 9, 9, 14, 15, 15, 21, 25, 26, 1, 1, 1, 1, 26, 25, 21, 14, 14, 14, 14, 18, 14, 17, 20, 19, 15, 16, 19, 20, 16, 14, 24, 26, 24, 12, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 10, 12, 25, 26, 23, 14, 21, 21, 20, 20, 21, 20, 20, 17, 14, 14, 18, 9, 9, 9, 14, 17, 21, 21, 21, 21, 17, 14, 9, 9, 9, 9, 9, 14, 20, 20, 20, 20, 16, 20, 21, 21, 14, 23, 26, 25, 12, 10, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 6, 12, 26, 1, 24, 14, 15, 19, 20, 20, 16, 15, 19, 19, 17, 17, 14, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 14, 14, 14, 20, 19, 15, 19, 19, 16, 16, 19, 21, 14, 21, 26, 26, 12, 6, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 1, 1, 23, 9, 15, 19, 15, 15, 15, 19, 20, 21, 21, 17, 14, 14, 14, 14, 14, 9, 14, 14, 14, 14, 14, 17, 20, 21, 21, 16, 16, 16, 19, 19, 19, 15, 14, 23, 26, 26, 7, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 24, 1, 1, 24, 14, 15, 16, 15, 15, 15, 16, 21, 21, 21, 19, 20, 20, 20, 20, 17, 17, 17, 17, 20, 20, 21, 21, 21, 20, 15, 19, 16, 16, 19, 20, 14, 23, 26, 1, 7, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 7, 7, 1, 1, 25, 17, 17, 16, 16, 15, 16, 20, 21, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 16, 16, 16, 16, 20, 14, 17, 25, 1, 1, 7, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 1, 27, 26, 23, 14, 17, 19, 16, 15, 20, 20, 20, 16, 16, 20, 20, 20, 20, 19, 19, 16, 16, 16, 16, 16, 19, 16, 20, 17, 14, 21, 26, 1, 26, 7, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 7, 26, 27, 1, 25, 17, 14, 15, 15, 16, 19, 19, 20, 16, 16, 20, 20, 20, 16, 16, 16, 16, 16, 16, 19, 16, 14, 17, 21, 25, 1, 27, 26, 7, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 12, 6, 27, 27, 26, 24, 15, 15, 15, 15, 15, 16, 16, 16, 19, 19, 19, 16, 16, 16, 16, 15, 15, 15, 15, 21, 24, 26, 27, 27, 6, 11, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 7, 1, 27, 27, 1, 25, 23, 15, 15, 15, 15, 15, 15, 15, 15, 17, 14, 14, 17, 17, 20, 23, 25, 1, 27, 27, 26, 7, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 11, 11, 1, 27, 28, 27, 1, 26, 25, 23, 21, 21, 20, 16, 19, 23, 23, 24, 26, 1, 27, 28, 27, 1, 11, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 11, 11, 10, 27, 28, 28, 28, 28, 27, 27, 27, 27, 27, 27, 27, 28, 28, 27, 27, 26, 11, 11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 7, 7, 11, 26, 1, 27, 27, 28, 28, 27, 27, 1, 1, 6, 11, 11, 6, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0),
		(0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 1, 2, 24, 24, 21, 23, 24, 24, 25, 26, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0)
	);
	
	signal cor_indice : integer := 0;
	type cor_int is array(0 to 2) of integer range 0 to 255;
	type matriz_cores is array(0 to N_CORES-1) of cor_int;
	constant obj_cores: matriz_cores :=
	(
		(0, 187, 204), --0
		(117, 177, 116),
		(88, 111, 87),
		(48, 81, 45),
		(7, 186, 202),--3
		(21, 182, 192),
		(37, 163, 155),
		(35, 141, 110),
		(27, 96, 24),
		(26, 109, 21),
		(30, 175, 179),
		(37, 151, 132),
		(29, 124, 86),
		(23, 83, 20),
		(32, 118, 28),
		(32, 131, 25),
		(36, 132, 30),
		(37, 122, 32),
		(33, 107, 29),
		(39, 134, 34),
		(38, 130, 33),
		(43, 130, 38),
		(17, 65, 14),
		(50, 138, 46),
		(60, 139, 57),
		(76, 152, 73),
		(97, 170, 95),
		(148, 201, 146),
		(181, 218, 181),
		(231, 245, 231)
	);

	
	signal pix_x: unsigned(9 downto 0) := unsigned( pixel_x );
	signal pix_y: unsigned(9 downto 0) := unsigned( pixel_y );
	
	begin				
		pix_x 	<= unsigned( pixel_x );
		pix_y 	<= unsigned( pixel_y );
		obj_Ymax <= obj_Ymin + LINHAS;
		obj_Xmax <= obj_Xmin + COLUNAS;
		
		forced_rst <= '1' when goal_tick = "10" else
						  '1'	when goal_tick = "01" else
						  '0';
		
		-- Atualizador de Registradores
		process( clk, reset, forced_rst, stop_game )
		begin
			if( reset = '1' or forced_rst = '1' or stop_game = '1' ) then
				obj_Ymin <= (480-LINHAS)/2;
				obj_Xmin <= 640 - 50 - COLUNAS;
				
			elsif( clk'event and clk='1' ) then
				obj_Ymin <= obj_Ymin_next;
				obj_Xmin <= obj_Xmin_next;
			end if;
		end process;
		
		-- Atualizador Posicao
		process( pad1_Rx_EN , pad1_Rx, pad1_Ry_EN, pad1_Ry,
					obj_Ymin, obj_Xmin, refresh_tick_pad )
		begin
			obj_Ymin_next <= obj_Ymin;
			obj_Xmin_next <= obj_Xmin;
			
			if( refresh_tick_pad = '1' ) then
				if( pad1_Rx_EN = '1' ) then
					if(     pad1_Rx = '0' ) then
						if( obj_Xmin < frontier_Xmax ) then obj_Xmin_next <= obj_Xmin + 1;
						else											obj_Xmin_next <= frontier_Xmax;
						end if;
					else
						if( obj_Xmin > frontier_Xmin ) then obj_Xmin_next <= obj_Xmin - 1;
						else											obj_Xmin_next <= frontier_Xmin;
						end if;
					end if;
				end if;
			
				if( pad1_Ry_EN = '1' ) then
					if(     pad1_Ry = '1' ) then
						if( obj_Ymin < frontier_Ymax ) then obj_Ymin_next <= obj_Ymin + 1;
						else											obj_Ymin_next <= frontier_Ymax;
						end if;
					else
						if( obj_Ymin > frontier_Ymin ) then obj_Ymin_next <= obj_Ymin - 1;
						else											obj_Ymin_next <= frontier_Ymin;
						end if;
					end if;
				end if;
			end if;
			
		end process;

		--Verifica saída de video
		process( pix_x, pix_y, cor_indice ,
				   obj_Xmin, obj_Xmax, obj_Ymin, obj_Ymax )
		begin
			obj_on		<= '0';
			obj_RGB(0)  <= "00000000";
			obj_RGB(1)  <= "00000000";
			obj_RGB(2)	<= "00000000";
			cor_indice	<= 0;
			
			if( (obj_Xmin <= pix_x) and (pix_x <= obj_Xmax) and
				 (obj_Ymin <= pix_y) and (pix_y <= obj_Ymax) ) then
				 
				cor_indice	<= obj_matriz( to_integer( pix_Y ) - obj_Ymin )
												 ( to_integer( pix_X ) - obj_Xmin );
												 
				case cor_indice is
					when 0  		=> obj_on <= '0';
					when 3 		=> obj_on <= '0';
					when others => obj_on <= '1';
				end case;
				
				obj_RGB(0) <= RGB_UNSIGNED( obj_cores(cor_indice)(0) );
				obj_RGB(1) <= RGB_UNSIGNED( obj_cores(cor_indice)(1) );
				obj_RGB(2) <= RGB_UNSIGNED( obj_cores(cor_indice)(2) );
				
			end if;
			
		end process;
		pad_Y <= std_logic_vector( to_unsigned( obj_Ymin , 10) );
		pad_X <= std_logic_vector( to_unsigned( obj_Xmin , 10) );
end arch;