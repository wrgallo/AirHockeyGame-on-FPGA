library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.TIPOS.all;

entity table is
	port(
		pixel_x, pixel_y:		 in std_logic_vector(9 downto 0);
		
		table_on:				out std_logic;
		table_RGB:				out TYPE_COR
	);
	
end table;

architecture arch of table is
	--Definicoes basicas da img
	constant LINHAS:  integer := 160;
   constant COLUNAS: integer := 240;
	constant N_CORES:	integer := 30;
	--Dimensoes da Imagem na tela
	constant Table_Ymin: integer := 26;
	constant Table_Ymax: integer := 26 + 428;
	constant Table_Xmin: integer := 0;
	constant Table_Xmax: integer := 0 + 640;
	--Definindo a img
	type linha_bitmap is array(0 to COLUNAS -1) of integer range 0 to N_CORES;
	type table_bitmap is array(0 to LINHAS  -1) of linha_bitmap;
	
   constant table_matriz: table_bitmap :=
	(
		(0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1),
		(0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1),
		(0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1),
		(0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1),
		(0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1),
		(0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1),
		(0, 1, 1, 1, 1, 1, 0, 3, 4, 5, 5, 6, 7, 5, 8, 4, 5, 6, 9, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 6, 5, 4, 6, 6, 4, 10, 4, 4, 6, 9, 4, 4, 6, 6, 4, 4, 4, 4, 4, 4, 8, 8, 10, 10, 4, 4, 6, 6, 10, 6, 6, 10, 10, 6, 9, 4, 10, 10, 4, 4, 10, 10, 3, 10, 4, 9, 4, 10, 3, 10, 10, 9, 9, 4, 4, 10, 4, 10, 4, 11, 9, 4, 10, 4, 5, 5, 5, 8, 3, 3, 4, 3, 10, 4, 9, 10, 4, 9, 4, 10, 4, 8, 8, 10, 10, 3, 3, 6, 10, 3, 5, 5, 10, 10, 4, 9, 10, 3, 3, 10, 10, 10, 10, 10, 3, 10, 4, 3, 4, 4, 4, 10, 3, 10, 4, 3, 3, 3, 3, 3, 3, 3, 10, 4, 6, 4, 10, 3, 3, 10, 10, 10, 4, 10, 10, 10, 10, 3, 10, 3, 3, 10, 4, 3, 3, 10, 3, 3, 10, 3, 3, 3, 4, 4, 10, 10, 4, 10, 4, 8, 3, 10, 10, 4, 5, 4, 6, 5, 10, 10, 10, 10, 4, 4, 4, 4, 4, 9, 10, 3, 10, 10, 3, 4, 10, 3, 10, 4, 4, 4, 6, 9, 10, 3, 10, 3, 10, 3, 3, 3, 10, 9, 3, 12, 0, 1, 1, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 12, 13, 14, 14, 14, 15, 15, 16, 17, 18, 14, 14, 14, 15, 14, 14, 14, 14, 14, 15, 14, 14, 14, 14, 14, 15, 14, 15, 15, 17, 17, 14, 14, 14, 14, 15, 14, 15, 14, 14, 14, 14, 17, 15, 14, 15, 17, 15, 17, 15, 14, 15, 17, 17, 14, 19, 15, 15, 14, 19, 14, 17, 19, 20, 20, 21, 17, 11, 17, 17, 17, 17, 13, 17, 13, 14, 15, 13, 15, 17, 17, 17, 15, 14, 14, 15, 15, 17, 15, 15, 17, 15, 13, 11, 17, 13, 19, 14, 14, 17, 17, 14, 15, 17, 11, 11, 11, 11, 11, 11, 15, 20, 22, 6, 11, 15, 14, 15, 15, 17, 17, 17, 17, 13, 11, 17, 17, 11, 17, 11, 13, 19, 18, 15, 17, 13, 15, 15, 17, 13, 22, 9, 11, 13, 17, 17, 17, 17, 17, 6, 11, 20, 23, 23, 9, 17, 19, 6, 11, 11, 17, 6, 6, 11, 11, 11, 4, 9, 6, 10, 24, 10, 5, 24, 8, 17, 19, 11, 4, 9, 9, 10, 9, 22, 10, 9, 16, 15, 13, 17, 14, 15, 23, 9, 24, 17, 11, 19, 11, 6, 17, 19, 13, 6, 11, 13, 10, 9, 20, 11, 11, 11, 14, 15, 13, 15, 17, 17, 11, 11, 7, 24, 24, 20, 21, 15, 16, 11, 12, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 15, 15, 14, 14, 14, 15, 15, 19, 19, 15, 14, 15, 15, 15, 15, 13, 19, 18, 18, 19, 15, 14, 15, 15, 15, 14, 15, 13, 19, 15, 14, 15, 15, 19, 19, 14, 19, 19, 15, 19, 19, 17, 19, 14, 14, 15, 15, 15, 14, 15, 19, 14, 19, 14, 14, 15, 19, 14, 19, 14, 14, 18, 23, 22, 20, 20, 18, 15, 19, 13, 14, 15, 15, 15, 16, 15, 21, 15, 15, 13, 15, 20, 14, 14, 21, 18, 14, 18, 21, 21, 21, 18, 15, 13, 17, 15, 19, 15, 15, 15, 15, 15, 16, 22, 24, 24, 23, 20, 14, 21, 24, 16, 8, 25, 4, 15, 11, 11, 19, 19, 15, 19, 19, 24, 16, 8, 22, 16, 17, 19, 21, 15, 15, 15, 18, 19, 13, 6, 19, 14, 19, 16, 21, 15, 14, 17, 15, 21, 20, 8, 8, 8, 8, 16, 8, 24, 22, 5, 22, 8, 9, 13, 13, 18, 23, 10, 4, 9, 9, 9, 9, 22, 17, 15, 13, 9, 22, 22, 22, 24, 8, 8, 23, 19, 15, 11, 24, 24, 23, 21, 13, 21, 23, 23, 11, 20, 24, 15, 21, 9, 23, 8, 8, 21, 18, 24, 9, 21, 21, 22, 21, 18, 15, 9, 18, 22, 18, 21, 13, 9, 24, 24, 11, 13, 15, 20, 15, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 4, 19, 19, 15, 19, 19, 15, 13, 17, 19, 15, 15, 17, 15, 14, 14, 13, 19, 15, 15, 15, 14, 14, 15, 15, 19, 15, 15, 13, 15, 17, 15, 19, 13, 11, 13, 19, 13, 17, 15, 17, 11, 13, 15, 15, 14, 14, 13, 15, 11, 17, 19, 19, 15, 14, 14, 15, 17, 14, 19, 15, 15, 19, 6, 6, 9, 19, 13, 17, 15, 15, 11, 15, 14, 17, 11, 19, 14, 17, 15, 15, 19, 13, 19, 14, 15, 15, 19, 11, 11, 11, 6, 13, 18, 14, 15, 15, 17, 14, 14, 17, 13, 19, 19, 20, 11, 11, 20, 15, 13, 8, 11, 14, 25, 26, 27, 15, 21, 22, 15, 19, 11, 6, 13, 18, 13, 21, 18, 11, 17, 15, 14, 15, 21, 9, 11, 18, 18, 19, 11, 15, 14, 6, 23, 14, 14, 17, 6, 20, 9, 8, 4, 9, 22, 8, 8, 8, 13, 6, 23, 6, 9, 4, 13, 21, 20, 24, 9, 4, 9, 21, 23, 11, 14, 15, 9, 9, 13, 20, 21, 24, 8, 22, 13, 18, 13, 23, 9, 9, 6, 13, 6, 23, 18, 11, 9, 9, 20, 13, 13, 6, 9, 8, 9, 9, 20, 19, 6, 13, 19, 20, 20, 20, 13, 11, 6, 15, 15, 17, 15, 17, 23, 23, 20, 9, 23, 18, 15, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 14, 15, 13, 6, 11, 13, 15, 17, 14, 14, 14, 15, 17, 14, 14, 17, 19, 19, 13, 15, 14, 17, 15, 14, 13, 15, 15, 13, 11, 19, 19, 19, 17, 13, 15, 17, 11, 19, 19, 17, 19, 15, 19, 13, 17, 15, 14, 11, 11, 13, 15, 19, 15, 15, 14, 15, 19, 15, 15, 17, 11, 13, 20, 11, 19, 14, 17, 13, 17, 15, 15, 19, 19, 14, 15, 13, 14, 15, 14, 14, 16, 11, 11, 14, 14, 15, 11, 11, 11, 23, 11, 21, 21, 14, 14, 15, 13, 13, 14, 13, 13, 19, 20, 6, 23, 13, 15, 13, 23, 18, 6, 18, 25, 26, 27, 15, 22, 11, 15, 13, 17, 15, 9, 21, 19, 18, 23, 11, 13, 15, 13, 13, 15, 13, 18, 21, 9, 23, 24, 8, 19, 9, 15, 17, 14, 17, 9, 20, 8, 8, 8, 21, 8, 10, 8, 9, 6, 11, 9, 23, 6, 11, 11, 23, 23, 23, 21, 20, 9, 9, 15, 14, 9, 23, 21, 9, 19, 15, 13, 11, 6, 18, 15, 23, 8, 23, 21, 23, 9, 20, 21, 6, 23, 20, 20, 13, 20, 6, 9, 18, 11, 6, 20, 8, 6, 21, 9, 20, 23, 21, 20, 20, 6, 18, 6, 17, 14, 14, 17, 6, 21, 21, 9, 13, 23, 19, 14, 4, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 6, 14, 21, 24, 24, 24, 13, 15, 19, 11, 13, 15, 14, 17, 15, 14, 15, 19, 13, 17, 14, 14, 19, 15, 14, 17, 15, 11, 17, 15, 19, 13, 17, 13, 13, 15, 11, 15, 15, 19, 14, 17, 11, 11, 17, 13, 15, 15, 13, 11, 13, 19, 14, 13, 17, 15, 14, 19, 19, 19, 19, 13, 13, 15, 13, 15, 13, 17, 13, 11, 13, 14, 15, 19, 15, 14, 14, 15, 14, 14, 15, 11, 11, 15, 15, 14, 18, 20, 13, 19, 19, 21, 21, 19, 11, 19, 14, 15, 13, 15, 15, 11, 13, 23, 23, 21, 14, 14, 21, 14, 22, 11, 15, 25, 26, 27, 14, 22, 11, 15, 19, 19, 13, 21, 13, 6, 8, 20, 11, 17, 15, 23, 23, 19, 21, 19, 11, 4, 9, 8, 8, 5, 14, 19, 4, 17, 11, 6, 20, 8, 9, 22, 8, 9, 9, 8, 9, 6, 11, 19, 9, 20, 15, 11, 21, 23, 23, 6, 23, 23, 15, 15, 6, 23, 8, 11, 19, 15, 21, 4, 6, 19, 15, 11, 8, 9, 9, 9, 13, 13, 13, 11, 9, 4, 11, 21, 9, 23, 18, 11, 23, 19, 20, 13, 8, 9, 19, 13, 23, 6, 6, 11, 9, 8, 19, 14, 15, 14, 15, 17, 6, 9, 23, 19, 11, 14, 14, 14, 5, 0, 1, 1, 1, 1),
		(2, 2, 2, 2, 1, 0, 4, 22, 22, 11, 11, 13, 21, 19, 18, 13, 11, 13, 15, 17, 15, 14, 14, 19, 17, 15, 15, 15, 13, 15, 14, 11, 17, 13, 17, 19, 11, 15, 14, 13, 17, 13, 13, 15, 13, 21, 18, 15, 17, 17, 11, 17, 15, 19, 14, 15, 17, 19, 15, 19, 13, 13, 14, 15, 15, 15, 13, 19, 13, 15, 14, 13, 13, 17, 17, 15, 15, 13, 13, 14, 14, 14, 14, 14, 15, 19, 14, 6, 15, 14, 15, 17, 14, 17, 13, 19, 19, 19, 19, 13, 13, 23, 19, 14, 15, 15, 15, 19, 6, 9, 17, 14, 14, 15, 15, 18, 18, 22, 19, 7, 28, 25, 15, 11, 23, 13, 15, 13, 17, 14, 23, 4, 23, 15, 14, 19, 24, 8, 10, 8, 22, 6, 20, 21, 13, 11, 23, 18, 14, 6, 13, 23, 22, 22, 8, 8, 19, 11, 6, 13, 9, 9, 9, 9, 23, 19, 19, 20, 19, 15, 13, 6, 11, 9, 9, 19, 11, 13, 20, 19, 13, 11, 15, 14, 6, 23, 21, 11, 13, 11, 6, 9, 4, 4, 11, 19, 20, 9, 9, 9, 9, 9, 24, 9, 24, 19, 9, 13, 15, 4, 8, 21, 15, 11, 8, 9, 9, 6, 13, 11, 11, 13, 14, 15, 15, 15, 20, 9, 23, 20, 9, 13, 14, 14, 29, 0, 1, 1, 1, 1),
		(2, 2, 2, 2, 2, 0, 10, 22, 21, 13, 21, 19, 19, 20, 13, 18, 15, 17, 15, 13, 11, 19, 17, 14, 14, 19, 15, 19, 13, 14, 17, 13, 14, 17, 13, 19, 11, 17, 17, 13, 14, 17, 19, 15, 18, 21, 13, 19, 13, 17, 19, 15, 13, 19, 15, 14, 15, 13, 15, 15, 11, 11, 17, 15, 15, 15, 17, 15, 17, 15, 15, 15, 17, 19, 15, 14, 15, 15, 19, 14, 14, 19, 13, 14, 19, 17, 15, 14, 13, 15, 19, 13, 14, 14, 13, 11, 13, 15, 19, 13, 13, 13, 13, 18, 15, 15, 14, 17, 13, 19, 19, 15, 14, 18, 13, 19, 19, 19, 13, 17, 14, 15, 19, 24, 8, 4, 14, 15, 14, 14, 15, 18, 20, 20, 13, 20, 23, 8, 8, 22, 21, 6, 9, 23, 13, 13, 18, 19, 13, 15, 15, 4, 8, 16, 9, 13, 13, 20, 20, 6, 13, 11, 23, 6, 11, 19, 19, 21, 11, 15, 21, 8, 6, 6, 13, 20, 9, 20, 13, 13, 13, 14, 14, 17, 11, 9, 4, 4, 13, 6, 9, 9, 6, 23, 9, 8, 9, 13, 19, 9, 9, 8, 8, 22, 9, 23, 20, 21, 21, 13, 20, 20, 23, 15, 9, 8, 8, 9, 20, 11, 9, 9, 15, 15, 17, 20, 18, 14, 20, 4, 4, 4, 15, 15, 4, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 15, 19, 18, 21, 19, 20, 13, 19, 15, 14, 15, 15, 11, 13, 15, 11, 17, 14, 15, 15, 14, 15, 19, 14, 14, 14, 15, 19, 15, 19, 19, 17, 15, 14, 15, 14, 15, 18, 19, 13, 18, 19, 13, 15, 11, 11, 13, 15, 14, 14, 17, 14, 15, 13, 13, 17, 15, 19, 15, 14, 15, 15, 15, 13, 15, 19, 14, 14, 15, 15, 15, 14, 14, 17, 13, 15, 14, 15, 14, 14, 14, 15, 15, 19, 11, 15, 14, 15, 13, 15, 19, 21, 20, 23, 19, 13, 6, 15, 14, 14, 14, 15, 15, 15, 19, 13, 21, 21, 13, 21, 19, 13, 13, 14, 16, 18, 24, 24, 13, 14, 14, 14, 15, 15, 21, 13, 21, 23, 9, 21, 11, 23, 13, 18, 13, 13, 23, 9, 11, 15, 13, 6, 14, 13, 18, 13, 14, 14, 19, 6, 9, 9, 6, 20, 20, 11, 23, 9, 19, 21, 23, 9, 23, 20, 11, 6, 13, 21, 20, 6, 20, 20, 23, 19, 15, 19, 20, 15, 4, 3, 20, 20, 9, 9, 6, 6, 9, 9, 9, 23, 6, 9, 22, 8, 10, 10, 24, 21, 9, 6, 18, 20, 18, 21, 8, 6, 13, 13, 23, 9, 23, 8, 8, 8, 9, 14, 17, 17, 6, 15, 18, 19, 20, 20, 9, 15, 17, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 13, 18, 21, 18, 20, 20, 21, 21, 13, 13, 17, 15, 13, 13, 15, 13, 11, 19, 14, 15, 14, 15, 15, 14, 14, 15, 15, 14, 19, 17, 19, 15, 14, 14, 14, 14, 15, 15, 15, 18, 21, 15, 15, 19, 17, 19, 13, 19, 15, 17, 14, 15, 19, 14, 13, 13, 14, 15, 15, 14, 14, 15, 17, 19, 17, 14, 14, 15, 15, 14, 14, 15, 19, 17, 19, 15, 14, 14, 14, 14, 14, 14, 15, 19, 19, 19, 15, 14, 15, 13, 20, 20, 11, 20, 21, 21, 19, 14, 14, 15, 14, 15, 15, 17, 13, 13, 20, 13, 20, 11, 6, 22, 7, 25, 25, 15, 17, 17, 15, 14, 17, 17, 13, 20, 14, 15, 15, 13, 23, 11, 11, 19, 17, 15, 13, 11, 6, 13, 19, 23, 6, 17, 15, 17, 11, 19, 14, 15, 17, 13, 23, 6, 9, 9, 8, 8, 8, 23, 21, 20, 6, 6, 6, 23, 15, 15, 20, 23, 11, 6, 23, 21, 21, 9, 21, 20, 9, 20, 15, 11, 13, 9, 11, 20, 11, 9, 23, 20, 23, 8, 4, 4, 8, 9, 24, 9, 9, 9, 6, 6, 15, 6, 11, 21, 21, 6, 11, 18, 23, 20, 23, 8, 4, 23, 18, 9, 17, 17, 13, 6, 21, 15, 20, 13, 19, 6, 18, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 4, 15, 13, 17, 13, 19, 18, 21, 13, 6, 11, 13, 15, 17, 13, 15, 17, 13, 15, 15, 14, 15, 19, 17, 14, 15, 15, 14, 15, 17, 11, 17, 14, 14, 14, 14, 19, 17, 19, 19, 19, 19, 14, 15, 21, 21, 13, 19, 19, 15, 15, 17, 15, 13, 15, 14, 14, 14, 14, 14, 14, 14, 14, 17, 17, 14, 14, 14, 13, 17, 14, 19, 17, 13, 19, 14, 14, 13, 15, 19, 14, 14, 15, 14, 19, 13, 11, 13, 14, 13, 6, 11, 20, 21, 15, 19, 19, 13, 15, 14, 14, 14, 15, 17, 17, 17, 13, 23, 20, 9, 16, 17, 14, 25, 26, 27, 14, 17, 17, 15, 19, 11, 8, 21, 19, 17, 19, 19, 18, 21, 18, 13, 20, 19, 19, 23, 11, 20, 18, 11, 23, 13, 15, 6, 14, 13, 14, 15, 19, 9, 6, 11, 20, 13, 11, 11, 23, 9, 9, 8, 4, 20, 19, 15, 14, 17, 20, 6, 9, 9, 11, 9, 18, 9, 23, 19, 23, 8, 4, 13, 15, 15, 13, 19, 23, 9, 9, 11, 24, 8, 9, 9, 4, 6, 9, 23, 20, 9, 8, 6, 15, 23, 13, 6, 6, 19, 21, 11, 21, 8, 8, 20, 11, 9, 9, 18, 9, 19, 17, 19, 20, 20, 13, 14, 15, 19, 9, 15, 4, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 4, 15, 15, 17, 13, 13, 13, 11, 20, 13, 11, 11, 19, 14, 17, 15, 17, 15, 19, 11, 14, 15, 13, 13, 15, 15, 15, 14, 19, 13, 13, 15, 14, 14, 14, 15, 19, 13, 13, 17, 13, 15, 15, 15, 21, 11, 21, 19, 13, 21, 15, 15, 15, 14, 17, 15, 17, 15, 14, 14, 14, 14, 14, 14, 14, 14, 19, 14, 15, 15, 19, 11, 17, 19, 14, 15, 17, 19, 13, 6, 13, 14, 15, 14, 19, 11, 6, 17, 15, 17, 11, 21, 18, 18, 19, 17, 13, 17, 14, 15, 11, 13, 14, 13, 17, 19, 13, 20, 19, 16, 15, 14, 15, 25, 26, 27, 14, 15, 14, 13, 6, 13, 8, 23, 14, 11, 19, 15, 20, 18, 14, 21, 20, 6, 13, 21, 23, 15, 19, 23, 11, 13, 20, 6, 17, 19, 15, 15, 19, 11, 23, 21, 23, 9, 6, 11, 13, 13, 24, 22, 9, 19, 15, 15, 15, 6, 11, 19, 6, 23, 8, 23, 13, 6, 14, 19, 8, 9, 20, 11, 15, 14, 11, 13, 6, 6, 23, 9, 4, 4, 4, 24, 24, 11, 22, 6, 9, 11, 6, 20, 13, 20, 20, 6, 9, 9, 13, 13, 21, 11, 8, 6, 13, 11, 20, 23, 11, 13, 13, 18, 13, 23, 6, 18, 15, 23, 22, 17, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 6, 14, 14, 15, 19, 13, 21, 13, 11, 11, 13, 17, 15, 15, 17, 15, 15, 17, 11, 13, 15, 19, 17, 19, 14, 15, 15, 15, 19, 15, 15, 15, 14, 14, 14, 15, 17, 19, 19, 13, 15, 15, 21, 21, 21, 19, 18, 20, 11, 21, 17, 15, 19, 15, 15, 19, 19, 13, 14, 14, 14, 14, 14, 14, 14, 15, 15, 15, 14, 15, 13, 15, 17, 15, 15, 17, 19, 13, 11, 13, 15, 15, 15, 14, 19, 15, 14, 19, 17, 14, 15, 15, 18, 21, 13, 17, 15, 14, 14, 11, 13, 13, 14, 15, 17, 15, 15, 14, 14, 19, 13, 5, 16, 25, 26, 27, 14, 15, 14, 21, 11, 19, 23, 18, 13, 15, 17, 15, 14, 11, 11, 13, 21, 20, 13, 19, 14, 21, 6, 20, 19, 15, 20, 11, 13, 15, 13, 23, 19, 15, 13, 20, 23, 9, 6, 6, 23, 23, 11, 16, 13, 15, 14, 15, 17, 6, 11, 20, 19, 9, 11, 11, 9, 15, 15, 9, 9, 9, 6, 14, 14, 19, 19, 23, 23, 21, 11, 9, 4, 8, 8, 8, 9, 6, 17, 23, 6, 23, 20, 19, 6, 20, 23, 23, 11, 9, 9, 20, 11, 21, 23, 23, 4, 4, 11, 23, 13, 13, 13, 19, 4, 11, 13, 8, 23, 9, 18, 13, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 9, 15, 18, 14, 14, 17, 13, 18, 19, 21, 15, 14, 14, 14, 14, 14, 15, 15, 17, 15, 15, 19, 14, 15, 14, 15, 14, 19, 19, 15, 17, 14, 14, 15, 19, 19, 17, 17, 17, 15, 15, 19, 19, 13, 15, 19, 20, 20, 19, 19, 19, 13, 13, 19, 15, 19, 19, 15, 14, 14, 14, 15, 14, 14, 15, 15, 14, 14, 14, 17, 15, 19, 17, 15, 13, 14, 19, 6, 6, 15, 14, 13, 11, 14, 14, 14, 15, 15, 19, 14, 14, 21, 21, 18, 19, 15, 14, 14, 11, 17, 15, 15, 19, 14, 14, 15, 17, 13, 13, 15, 13, 11, 14, 5, 28, 25, 14, 17, 17, 13, 13, 15, 18, 21, 13, 15, 14, 11, 13, 13, 6, 20, 13, 23, 11, 14, 21, 20, 21, 15, 21, 21, 13, 15, 11, 19, 15, 11, 11, 15, 23, 23, 20, 11, 4, 23, 20, 9, 6, 22, 6, 13, 15, 17, 15, 19, 11, 6, 6, 19, 11, 13, 13, 14, 13, 23, 11, 21, 15, 13, 17, 6, 11, 20, 13, 4, 9, 22, 21, 13, 22, 24, 24, 6, 11, 6, 6, 23, 11, 21, 21, 11, 9, 20, 11, 8, 4, 8, 21, 21, 23, 23, 9, 6, 21, 23, 19, 19, 11, 11, 11, 11, 19, 9, 11, 9, 18, 15, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 17, 16, 19, 14, 14, 11, 6, 13, 15, 18, 13, 15, 14, 15, 14, 14, 17, 15, 14, 15, 17, 15, 14, 14, 15, 15, 15, 14, 19, 13, 14, 14, 15, 15, 15, 15, 15, 15, 14, 15, 17, 21, 21, 15, 18, 13, 20, 21, 19, 15, 17, 17, 14, 17, 15, 17, 14, 17, 14, 15, 14, 14, 11, 13, 14, 14, 13, 11, 14, 14, 13, 15, 19, 18, 11, 13, 21, 15, 13, 20, 19, 17, 17, 14, 14, 14, 19, 17, 13, 14, 17, 17, 19, 13, 19, 15, 15, 17, 14, 15, 14, 19, 19, 13, 15, 17, 14, 17, 11, 15, 14, 11, 24, 18, 14, 14, 11, 23, 21, 21, 15, 18, 21, 23, 11, 11, 13, 6, 21, 18, 16, 24, 8, 22, 15, 21, 15, 15, 15, 13, 11, 15, 19, 6, 14, 15, 20, 23, 19, 13, 9, 6, 21, 18, 20, 4, 8, 23, 20, 20, 13, 11, 19, 11, 13, 8, 8, 23, 17, 17, 21, 6, 14, 23, 8, 23, 9, 13, 9, 13, 6, 19, 22, 8, 9, 9, 8, 10, 8, 22, 19, 19, 20, 16, 23, 23, 23, 21, 20, 11, 19, 13, 9, 9, 23, 10, 4, 11, 14, 23, 9, 13, 15, 15, 19, 18, 23, 21, 17, 14, 9, 8, 23, 20, 21, 15, 6, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 13, 16, 6, 13, 15, 14, 13, 17, 17, 21, 20, 20, 21, 15, 15, 14, 13, 13, 15, 17, 17, 19, 15, 14, 14, 14, 15, 15, 15, 15, 14, 13, 19, 17, 15, 15, 17, 15, 17, 13, 11, 13, 18, 20, 21, 13, 13, 20, 13, 11, 19, 14, 14, 15, 19, 14, 15, 19, 15, 14, 14, 15, 13, 19, 19, 14, 19, 13, 15, 17, 17, 14, 15, 20, 13, 21, 19, 21, 23, 9, 6, 19, 14, 14, 14, 19, 13, 6, 11, 14, 15, 6, 6, 15, 15, 14, 19, 15, 13, 13, 13, 15, 14, 15, 19, 14, 15, 14, 14, 22, 4, 6, 16, 15, 16, 15, 24, 24, 13, 21, 15, 20, 6, 20, 21, 23, 13, 15, 23, 19, 21, 4, 13, 15, 15, 19, 20, 13, 13, 15, 14, 18, 11, 13, 18, 19, 20, 8, 9, 20, 11, 8, 9, 20, 8, 9, 20, 23, 11, 6, 20, 23, 23, 23, 6, 23, 9, 23, 23, 15, 11, 23, 15, 23, 21, 23, 20, 9, 10, 21, 6, 3, 8, 22, 8, 22, 8, 10, 9, 24, 11, 19, 21, 11, 13, 9, 13, 18, 21, 6, 4, 6, 20, 23, 21, 13, 21, 13, 21, 14, 23, 20, 18, 19, 15, 23, 8, 8, 6, 15, 11, 8, 19, 13, 15, 22, 4, 3, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 11, 16, 20, 23, 11, 17, 14, 14, 13, 11, 11, 11, 20, 15, 19, 17, 13, 17, 17, 11, 11, 13, 17, 14, 14, 13, 13, 19, 19, 15, 14, 13, 13, 13, 13, 17, 15, 19, 17, 11, 17, 19, 23, 23, 20, 11, 20, 23, 23, 11, 17, 13, 15, 14, 15, 15, 15, 15, 14, 14, 15, 14, 15, 19, 17, 15, 14, 15, 6, 17, 14, 13, 9, 11, 13, 21, 13, 23, 21, 21, 13, 19, 11, 11, 19, 6, 11, 13, 19, 14, 14, 13, 15, 19, 13, 19, 13, 19, 11, 20, 6, 15, 14, 15, 19, 14, 14, 17, 13, 22, 6, 16, 6, 25, 29, 15, 20, 20, 11, 9, 23, 13, 23, 19, 13, 11, 9, 20, 20, 19, 17, 15, 14, 6, 13, 20, 15, 18, 21, 15, 18, 21, 20, 19, 20, 6, 21, 11, 11, 23, 11, 11, 6, 4, 23, 9, 20, 15, 9, 9, 6, 23, 9, 13, 9, 19, 13, 20, 8, 8, 6, 21, 23, 9, 4, 23, 11, 11, 13, 19, 9, 10, 3, 8, 24, 10, 9, 22, 9, 24, 19, 21, 9, 11, 13, 11, 13, 13, 6, 20, 6, 9, 23, 18, 14, 14, 13, 6, 8, 19, 19, 13, 21, 11, 13, 20, 23, 8, 23, 6, 15, 13, 18, 13, 13, 22, 6, 3, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 8, 17, 21, 19, 13, 13, 17, 15, 15, 15, 19, 13, 20, 6, 15, 6, 13, 11, 13, 13, 23, 21, 15, 15, 14, 19, 15, 19, 13, 17, 15, 15, 19, 11, 6, 6, 11, 13, 13, 13, 17, 13, 13, 21, 11, 21, 15, 13, 11, 13, 19, 15, 17, 19, 14, 14, 15, 14, 14, 14, 19, 14, 14, 15, 13, 19, 17, 11, 13, 15, 14, 15, 17, 6, 20, 9, 20, 20, 23, 11, 13, 18, 15, 11, 8, 11, 15, 19, 14, 14, 17, 14, 14, 13, 6, 11, 13, 13, 16, 22, 22, 22, 11, 13, 14, 14, 15, 13, 17, 11, 5, 19, 16, 25, 26, 27, 14, 16, 11, 11, 6, 11, 18, 20, 13, 8, 9, 23, 23, 19, 15, 15, 14, 17, 6, 23, 15, 19, 6, 21, 6, 23, 9, 11, 21, 13, 20, 18, 23, 4, 9, 11, 13, 23, 4, 11, 17, 11, 6, 11, 18, 21, 11, 6, 11, 21, 11, 14, 9, 8, 8, 11, 14, 8, 8, 8, 8, 9, 11, 9, 20, 13, 20, 8, 10, 22, 22, 8, 9, 22, 22, 21, 11, 23, 11, 11, 14, 15, 13, 6, 8, 8, 8, 4, 23, 23, 18, 14, 19, 21, 15, 14, 18, 13, 9, 6, 9, 9, 18, 23, 8, 13, 15, 11, 19, 20, 9, 9, 8, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 4, 17, 11, 17, 15, 17, 15, 20, 11, 21, 19, 15, 15, 13, 17, 4, 15, 13, 23, 18, 13, 19, 13, 21, 14, 13, 15, 18, 13, 20, 18, 13, 13, 19, 18, 19, 21, 20, 13, 13, 19, 13, 11, 20, 11, 20, 13, 13, 20, 21, 19, 15, 13, 19, 14, 14, 15, 14, 14, 14, 14, 17, 14, 15, 11, 24, 11, 11, 11, 14, 14, 11, 15, 15, 20, 21, 18, 20, 9, 6, 20, 6, 15, 17, 11, 17, 14, 15, 15, 15, 11, 13, 14, 17, 11, 19, 20, 9, 23, 11, 13, 20, 13, 14, 14, 13, 9, 9, 23, 11, 17, 17, 15, 25, 26, 27, 14, 15, 17, 23, 9, 9, 13, 6, 20, 23, 9, 9, 23, 21, 14, 14, 13, 11, 13, 23, 18, 9, 13, 6, 4, 23, 8, 6, 17, 19, 4, 11, 20, 6, 4, 20, 9, 23, 20, 6, 23, 8, 9, 23, 21, 11, 21, 20, 20, 15, 19, 23, 13, 6, 20, 15, 13, 9, 13, 6, 20, 22, 8, 6, 8, 9, 23, 6, 19, 13, 15, 21, 20, 20, 15, 6, 4, 20, 9, 8, 19, 9, 6, 11, 11, 23, 20, 19, 11, 6, 9, 13, 19, 9, 14, 15, 14, 19, 11, 13, 6, 13, 9, 8, 6, 17, 15, 6, 13, 21, 9, 13, 3, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 17, 15, 13, 19, 13, 19, 13, 23, 23, 17, 15, 13, 19, 15, 17, 15, 11, 13, 18, 15, 13, 23, 19, 14, 21, 11, 15, 18, 13, 13, 21, 13, 20, 21, 14, 19, 11, 20, 19, 11, 23, 20, 20, 13, 19, 19, 15, 21, 11, 20, 11, 21, 14, 14, 13, 14, 14, 15, 14, 15, 14, 14, 15, 9, 22, 6, 6, 14, 17, 15, 14, 17, 14, 18, 19, 23, 13, 11, 18, 13, 21, 14, 14, 14, 13, 13, 15, 6, 15, 14, 24, 11, 17, 13, 19, 9, 8, 20, 15, 13, 13, 14, 17, 13, 11, 9, 24, 4, 6, 17, 6, 14, 29, 26, 27, 14, 24, 23, 6, 9, 6, 11, 11, 8, 9, 9, 11, 20, 15, 14, 15, 11, 9, 9, 18, 15, 20, 11, 9, 13, 23, 20, 20, 23, 9, 13, 11, 23, 8, 9, 11, 20, 11, 13, 9, 10, 23, 13, 20, 13, 8, 8, 20, 18, 13, 20, 9, 21, 19, 13, 15, 13, 23, 14, 19, 21, 24, 8, 11, 8, 6, 13, 8, 6, 9, 23, 19, 19, 14, 21, 19, 19, 9, 8, 11, 11, 23, 9, 9, 9, 20, 13, 20, 23, 6, 6, 9, 19, 14, 19, 13, 19, 17, 14, 13, 19, 20, 9, 23, 19, 15, 19, 14, 6, 13, 19, 17, 3, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 13, 6, 19, 14, 15, 13, 23, 23, 20, 11, 15, 15, 17, 17, 14, 14, 11, 19, 18, 20, 19, 13, 19, 15, 20, 6, 20, 14, 18, 23, 21, 13, 13, 15, 19, 19, 18, 19, 11, 20, 11, 6, 21, 15, 18, 13, 21, 13, 20, 19, 15, 15, 20, 13, 19, 15, 14, 14, 17, 14, 17, 17, 15, 13, 21, 11, 19, 14, 13, 13, 15, 15, 11, 14, 19, 6, 13, 14, 14, 18, 14, 14, 13, 11, 6, 13, 19, 11, 11, 9, 19, 14, 15, 15, 17, 13, 20, 18, 11, 18, 15, 9, 8, 11, 19, 8, 10, 9, 6, 6, 19, 14, 7, 25, 25, 19, 24, 20, 23, 11, 6, 6, 11, 8, 23, 21, 21, 20, 19, 11, 6, 13, 24, 8, 11, 15, 14, 11, 11, 18, 11, 20, 23, 20, 9, 8, 9, 11, 8, 18, 6, 15, 23, 4, 6, 9, 9, 11, 23, 6, 4, 11, 14, 21, 23, 19, 14, 19, 15, 15, 18, 13, 21, 11, 17, 4, 10, 10, 6, 4, 9, 20, 8, 8, 20, 23, 20, 14, 11, 15, 19, 13, 13, 13, 18, 6, 11, 9, 8, 23, 20, 9, 9, 19, 13, 9, 20, 23, 20, 14, 14, 15, 11, 15, 17, 19, 20, 20, 23, 19, 11, 13, 14, 15, 17, 19, 17, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 4, 13, 13, 19, 13, 14, 15, 18, 18, 21, 17, 13, 14, 15, 11, 13, 15, 15, 15, 18, 11, 20, 15, 11, 13, 11, 23, 20, 13, 14, 21, 19, 11, 19, 13, 20, 11, 19, 21, 13, 13, 21, 19, 15, 18, 20, 11, 18, 18, 13, 11, 18, 13, 6, 14, 14, 19, 11, 15, 14, 15, 15, 17, 15, 19, 15, 14, 14, 14, 19, 11, 11, 13, 19, 17, 14, 14, 14, 13, 21, 21, 11, 19, 23, 6, 20, 18, 14, 14, 9, 9, 24, 15, 14, 15, 6, 19, 14, 15, 19, 21, 9, 4, 9, 8, 16, 8, 24, 20, 6, 13, 17, 17, 5, 16, 16, 17, 17, 11, 20, 11, 6, 11, 15, 23, 9, 8, 9, 15, 20, 9, 8, 8, 22, 22, 6, 15, 14, 19, 20, 6, 9, 21, 23, 23, 4, 8, 9, 11, 18, 21, 20, 21, 6, 4, 11, 13, 6, 20, 15, 6, 19, 14, 23, 9, 23, 9, 19, 23, 18, 15, 6, 11, 6, 9, 11, 23, 8, 8, 11, 11, 23, 23, 23, 8, 23, 9, 21, 19, 21, 6, 23, 11, 6, 18, 19, 6, 21, 18, 13, 20, 6, 23, 6, 9, 6, 19, 19, 23, 11, 14, 15, 14, 6, 11, 15, 11, 13, 20, 18, 19, 11, 13, 15, 15, 15, 22, 17, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 17, 15, 15, 17, 15, 15, 13, 14, 15, 17, 13, 11, 13, 15, 15, 17, 13, 21, 15, 18, 11, 13, 11, 17, 11, 13, 11, 13, 13, 19, 17, 19, 17, 20, 20, 13, 23, 9, 23, 19, 17, 15, 15, 21, 13, 20, 13, 21, 13, 21, 6, 6, 15, 14, 19, 11, 19, 14, 14, 11, 17, 14, 14, 14, 15, 14, 17, 17, 17, 11, 11, 17, 14, 14, 17, 15, 17, 19, 13, 6, 6, 20, 6, 4, 6, 22, 22, 15, 17, 23, 9, 11, 14, 14, 17, 6, 11, 14, 14, 11, 9, 8, 9, 9, 6, 15, 18, 9, 8, 11, 19, 4, 16, 18, 16, 17, 15, 6, 11, 11, 11, 13, 14, 20, 8, 10, 19, 13, 10, 24, 9, 8, 6, 14, 14, 18, 23, 9, 13, 8, 20, 23, 9, 8, 4, 9, 6, 21, 15, 15, 15, 6, 13, 11, 22, 24, 11, 11, 6, 23, 19, 4, 10, 8, 9, 10, 8, 23, 20, 15, 15, 23, 4, 9, 20, 20, 13, 9, 13, 9, 9, 6, 21, 9, 4, 21, 13, 6, 23, 9, 4, 20, 21, 20, 9, 23, 23, 13, 13, 20, 21, 21, 9, 11, 21, 23, 23, 13, 15, 13, 15, 17, 15, 15, 11, 21, 23, 9, 20, 6, 18, 21, 21, 15, 13, 16, 11, 3, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 4, 13, 13, 13, 15, 15, 14, 15, 13, 11, 15, 19, 13, 19, 17, 14, 17, 13, 19, 9, 23, 15, 13, 19, 19, 19, 11, 11, 21, 6, 11, 14, 13, 6, 11, 19, 6, 9, 23, 20, 13, 15, 15, 20, 9, 11, 21, 19, 11, 14, 15, 13, 14, 14, 17, 15, 15, 15, 19, 13, 13, 11, 15, 14, 14, 14, 13, 13, 19, 15, 14, 15, 15, 6, 15, 14, 17, 13, 18, 23, 9, 4, 23, 4, 6, 21, 22, 8, 22, 15, 20, 23, 19, 14, 14, 13, 17, 19, 17, 17, 19, 16, 20, 13, 15, 15, 14, 8, 8, 8, 18, 22, 23, 29, 28, 25, 17, 16, 16, 19, 23, 8, 4, 6, 9, 21, 18, 15, 4, 10, 4, 19, 20, 18, 19, 21, 9, 11, 20, 13, 13, 20, 9, 19, 21, 18, 20, 13, 18, 15, 6, 9, 11, 11, 4, 10, 10, 4, 19, 6, 19, 9, 8, 24, 8, 10, 10, 10, 23, 21, 6, 14, 21, 19, 20, 11, 9, 8, 6, 23, 9, 20, 20, 18, 9, 13, 13, 4, 9, 9, 20, 6, 11, 23, 19, 23, 6, 20, 11, 6, 9, 9, 23, 13, 15, 15, 13, 13, 13, 21, 23, 13, 19, 14, 11, 9, 9, 13, 21, 13, 20, 23, 9, 23, 21, 20, 24, 11, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 6, 8, 4, 23, 23, 11, 19, 17, 13, 15, 14, 14, 14, 13, 17, 19, 17, 13, 23, 20, 19, 11, 19, 14, 17, 9, 20, 13, 11, 13, 14, 13, 6, 21, 13, 21, 20, 23, 23, 9, 11, 19, 21, 21, 6, 23, 11, 21, 18, 19, 14, 14, 19, 17, 15, 19, 19, 17, 13, 15, 19, 17, 14, 14, 14, 19, 15, 20, 23, 6, 13, 20, 20, 15, 13, 21, 20, 9, 19, 20, 6, 23, 11, 19, 9, 24, 8, 9, 17, 15, 15, 13, 13, 15, 14, 17, 9, 19, 13, 11, 15, 18, 11, 15, 18, 19, 19, 23, 18, 19, 8, 16, 25, 26, 27, 14, 20, 13, 22, 22, 10, 10, 23, 8, 6, 17, 17, 17, 19, 16, 6, 11, 19, 6, 15, 15, 13, 21, 20, 18, 20, 11, 19, 9, 6, 6, 18, 21, 6, 9, 4, 23, 23, 9, 3, 10, 9, 15, 21, 10, 11, 19, 8, 10, 8, 8, 8, 19, 14, 13, 23, 20, 11, 6, 11, 6, 10, 23, 19, 20, 23, 6, 19, 19, 18, 9, 6, 9, 6, 9, 15, 9, 23, 20, 20, 23, 9, 20, 13, 9, 9, 13, 19, 13, 9, 6, 19, 18, 18, 13, 13, 17, 14, 11, 9, 6, 19, 18, 9, 9, 9, 23, 23, 11, 6, 24, 17, 8, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 4, 11, 24, 21, 20, 23, 11, 13, 13, 13, 15, 15, 14, 15, 17, 14, 15, 15, 17, 20, 13, 13, 11, 13, 13, 14, 18, 21, 6, 11, 15, 13, 17, 15, 19, 13, 11, 6, 23, 23, 13, 13, 13, 13, 19, 21, 6, 20, 19, 11, 14, 19, 17, 19, 19, 14, 15, 14, 14, 19, 19, 14, 15, 15, 14, 15, 23, 9, 8, 9, 23, 23, 20, 18, 20, 20, 18, 20, 20, 9, 21, 21, 15, 15, 9, 4, 8, 8, 23, 17, 18, 21, 21, 15, 6, 14, 14, 19, 19, 15, 11, 24, 21, 14, 18, 6, 6, 13, 11, 17, 11, 20, 16, 25, 26, 27, 14, 16, 11, 8, 8, 24, 8, 9, 18, 14, 15, 17, 13, 13, 6, 18, 19, 20, 19, 23, 20, 15, 11, 23, 18, 21, 20, 23, 8, 9, 18, 18, 6, 8, 20, 9, 23, 8, 21, 8, 10, 19, 19, 9, 6, 9, 20, 24, 9, 24, 22, 16, 16, 13, 11, 4, 11, 20, 4, 4, 21, 11, 11, 20, 23, 23, 20, 18, 18, 6, 9, 9, 9, 9, 6, 23, 11, 13, 4, 4, 6, 20, 6, 11, 13, 21, 6, 9, 9, 9, 23, 20, 20, 19, 19, 6, 15, 15, 19, 19, 20, 21, 18, 21, 6, 6, 6, 11, 23, 18, 22, 17, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 17, 19, 21, 23, 23, 11, 11, 15, 15, 21, 20, 21, 16, 13, 19, 14, 14, 14, 15, 15, 17, 15, 14, 17, 17, 15, 14, 19, 17, 17, 11, 13, 15, 11, 11, 11, 13, 11, 6, 18, 20, 11, 19, 21, 18, 14, 15, 15, 14, 14, 15, 13, 13, 15, 15, 14, 15, 13, 19, 14, 14, 15, 15, 14, 14, 16, 9, 9, 24, 21, 20, 11, 6, 9, 9, 11, 18, 15, 13, 9, 19, 14, 22, 8, 8, 9, 9, 9, 22, 16, 13, 21, 21, 15, 14, 14, 19, 15, 13, 23, 13, 14, 18, 15, 19, 9, 20, 18, 9, 5, 19, 16, 25, 26, 27, 14, 16, 17, 23, 20, 19, 15, 14, 14, 13, 9, 8, 10, 8, 21, 15, 9, 6, 19, 21, 20, 14, 13, 11, 6, 9, 20, 23, 4, 19, 16, 8, 9, 8, 24, 23, 4, 23, 8, 23, 13, 15, 23, 11, 13, 20, 23, 21, 9, 9, 4, 11, 6, 20, 22, 6, 22, 19, 22, 9, 20, 20, 21, 11, 13, 13, 23, 22, 21, 8, 8, 6, 9, 4, 9, 10, 16, 9, 10, 8, 8, 9, 22, 13, 17, 13, 4, 8, 9, 9, 20, 11, 6, 20, 13, 17, 11, 13, 17, 11, 15, 18, 19, 15, 19, 9, 9, 9, 6, 11, 19, 19, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 8, 17, 16, 21, 20, 20, 11, 6, 17, 17, 9, 13, 20, 23, 22, 6, 17, 14, 13, 15, 17, 11, 17, 15, 14, 14, 19, 15, 14, 14, 14, 15, 13, 13, 15, 17, 17, 17, 21, 15, 15, 21, 18, 15, 21, 13, 17, 17, 14, 17, 13, 15, 11, 17, 11, 19, 19, 17, 19, 15, 17, 9, 13, 15, 14, 14, 14, 20, 11, 19, 15, 13, 6, 23, 6, 9, 8, 11, 19, 19, 19, 14, 17, 9, 13, 13, 23, 8, 18, 18, 15, 21, 15, 15, 19, 19, 15, 15, 13, 14, 23, 19, 11, 21, 13, 19, 15, 14, 14, 11, 5, 11, 16, 6, 25, 25, 15, 6, 19, 18, 18, 18, 19, 15, 19, 9, 9, 8, 8, 22, 18, 19, 11, 21, 11, 20, 18, 19, 14, 13, 4, 9, 6, 23, 15, 13, 8, 8, 8, 8, 8, 23, 8, 8, 23, 15, 14, 15, 21, 6, 9, 13, 23, 11, 21, 9, 11, 17, 13, 22, 24, 22, 9, 6, 11, 9, 23, 20, 6, 9, 21, 19, 19, 24, 24, 8, 8, 4, 9, 23, 8, 9, 8, 8, 8, 10, 8, 8, 24, 11, 11, 9, 20, 9, 8, 23, 21, 20, 8, 13, 15, 21, 15, 9, 23, 18, 13, 13, 20, 23, 18, 18, 23, 23, 20, 18, 16, 11, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 4, 17, 14, 21, 23, 9, 22, 16, 22, 16, 11, 20, 23, 23, 20, 13, 17, 17, 4, 17, 19, 15, 14, 17, 13, 17, 13, 17, 14, 13, 14, 14, 15, 17, 15, 14, 15, 13, 13, 21, 11, 19, 19, 16, 18, 18, 15, 14, 14, 14, 14, 15, 14, 15, 17, 14, 13, 19, 15, 13, 11, 13, 15, 11, 14, 14, 17, 19, 17, 17, 13, 13, 13, 13, 20, 23, 13, 20, 11, 15, 14, 14, 15, 15, 11, 6, 17, 14, 14, 19, 21, 18, 15, 15, 11, 17, 19, 14, 13, 15, 15, 20, 23, 13, 18, 15, 14, 14, 14, 11, 5, 19, 13, 5, 16, 16, 17, 6, 11, 15, 18, 19, 21, 11, 19, 19, 9, 9, 11, 13, 11, 23, 20, 15, 19, 23, 9, 23, 15, 19, 23, 6, 19, 19, 19, 6, 9, 24, 10, 10, 10, 11, 23, 9, 18, 14, 18, 18, 11, 20, 23, 6, 18, 11, 23, 11, 21, 13, 9, 8, 10, 22, 10, 4, 24, 13, 9, 11, 9, 9, 6, 4, 19, 9, 24, 8, 10, 4, 11, 13, 11, 9, 10, 10, 24, 9, 6, 22, 9, 8, 23, 20, 8, 9, 15, 20, 23, 6, 11, 15, 19, 23, 23, 23, 23, 19, 11, 9, 21, 8, 9, 21, 15, 15, 13, 19, 24, 4, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 11, 11, 13, 15, 19, 24, 8, 24, 8, 15, 18, 19, 13, 11, 13, 14, 14, 19, 19, 23, 13, 14, 14, 14, 14, 14, 15, 13, 15, 15, 17, 19, 14, 14, 15, 14, 13, 19, 15, 21, 19, 13, 13, 15, 14, 14, 14, 14, 17, 15, 14, 15, 13, 17, 13, 14, 15, 13, 13, 13, 15, 19, 13, 14, 14, 14, 14, 15, 17, 13, 20, 20, 20, 20, 19, 13, 21, 15, 14, 14, 14, 17, 6, 17, 15, 14, 14, 17, 11, 6, 18, 21, 19, 20, 11, 11, 13, 14, 15, 23, 18, 20, 13, 21, 18, 15, 17, 17, 14, 19, 19, 11, 22, 14, 14, 17, 19, 21, 6, 6, 15, 20, 23, 19, 14, 13, 6, 5, 6, 6, 19, 13, 23, 6, 13, 13, 20, 13, 11, 11, 9, 19, 19, 9, 11, 20, 24, 24, 24, 24, 11, 17, 13, 15, 21, 15, 8, 6, 6, 8, 6, 9, 23, 4, 11, 18, 4, 8, 8, 8, 8, 24, 24, 9, 11, 6, 11, 20, 11, 9, 20, 4, 4, 9, 24, 8, 6, 20, 8, 23, 16, 9, 8, 8, 17, 19, 6, 4, 8, 8, 9, 23, 13, 13, 17, 6, 13, 19, 14, 9, 20, 9, 4, 21, 19, 11, 9, 23, 23, 6, 20, 18, 21, 13, 21, 22, 6, 3, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 19, 22, 21, 20, 13, 11, 11, 11, 11, 13, 17, 19, 19, 18, 15, 15, 14, 18, 13, 21, 18, 21, 16, 13, 14, 15, 13, 13, 15, 15, 13, 13, 13, 13, 19, 14, 14, 19, 15, 15, 15, 19, 14, 14, 14, 14, 15, 14, 14, 15, 13, 15, 19, 17, 15, 19, 13, 13, 13, 13, 19, 23, 22, 17, 14, 15, 14, 15, 6, 24, 22, 22, 21, 20, 13, 13, 19, 19, 14, 15, 14, 15, 17, 14, 14, 14, 17, 13, 13, 11, 20, 13, 11, 19, 21, 23, 23, 14, 15, 13, 22, 21, 11, 9, 13, 21, 21, 15, 14, 14, 17, 21, 4, 28, 25, 18, 22, 6, 13, 17, 15, 18, 23, 20, 20, 21, 15, 13, 9, 6, 19, 9, 8, 8, 4, 20, 18, 23, 4, 13, 14, 19, 6, 20, 18, 19, 15, 20, 23, 10, 5, 15, 17, 4, 9, 16, 10, 10, 24, 8, 24, 9, 4, 8, 13, 16, 8, 8, 10, 8, 8, 21, 22, 8, 8, 22, 19, 6, 9, 13, 23, 9, 8, 8, 9, 13, 15, 11, 6, 13, 19, 13, 6, 11, 15, 19, 8, 4, 4, 4, 9, 20, 11, 6, 15, 13, 20, 15, 19, 6, 13, 4, 9, 20, 11, 19, 13, 11, 9, 11, 23, 11, 19, 20, 20, 18, 17, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 17, 16, 19, 11, 23, 13, 17, 15, 14, 14, 14, 14, 13, 6, 11, 13, 14, 19, 6, 21, 23, 23, 9, 11, 14, 13, 19, 19, 13, 15, 17, 13, 11, 6, 11, 13, 14, 14, 17, 11, 11, 15, 14, 14, 15, 15, 17, 15, 15, 15, 13, 15, 14, 14, 15, 15, 15, 21, 11, 15, 13, 22, 19, 13, 19, 14, 14, 13, 13, 11, 23, 23, 11, 6, 11, 15, 19, 17, 15, 13, 14, 14, 14, 17, 17, 17, 15, 15, 19, 15, 15, 13, 11, 19, 21, 20, 15, 15, 17, 13, 22, 6, 13, 13, 19, 16, 23, 6, 14, 14, 14, 14, 25, 26, 27, 14, 9, 6, 15, 15, 13, 13, 19, 21, 21, 6, 9, 13, 23, 6, 13, 23, 24, 24, 9, 20, 20, 21, 14, 18, 14, 18, 8, 8, 9, 10, 9, 21, 6, 19, 14, 19, 11, 4, 23, 21, 8, 10, 4, 9, 8, 9, 9, 6, 14, 4, 8, 8, 8, 22, 22, 9, 22, 10, 8, 22, 14, 4, 13, 11, 11, 23, 8, 8, 18, 19, 11, 11, 17, 19, 11, 20, 18, 18, 6, 23, 20, 9, 9, 6, 20, 13, 23, 18, 15, 11, 18, 14, 20, 11, 18, 6, 20, 23, 23, 23, 20, 18, 9, 20, 19, 6, 11, 14, 23, 22, 6, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 11, 24, 19, 14, 14, 14, 14, 14, 14, 11, 13, 17, 6, 22, 11, 11, 15, 6, 19, 13, 13, 21, 8, 17, 17, 11, 17, 19, 19, 14, 17, 13, 13, 19, 15, 13, 13, 14, 15, 15, 15, 14, 14, 13, 6, 23, 20, 13, 23, 6, 17, 14, 14, 14, 14, 14, 19, 13, 14, 19, 18, 18, 18, 17, 15, 14, 14, 14, 13, 15, 17, 11, 11, 17, 14, 17, 17, 17, 11, 13, 14, 15, 11, 11, 17, 9, 18, 13, 9, 18, 14, 15, 14, 23, 15, 19, 23, 17, 17, 9, 22, 13, 15, 14, 15, 9, 24, 11, 15, 19, 6, 14, 29, 26, 27, 14, 22, 15, 15, 17, 11, 13, 13, 13, 15, 6, 20, 23, 21, 13, 13, 6, 21, 21, 14, 14, 20, 13, 19, 6, 18, 6, 24, 10, 10, 8, 4, 6, 14, 19, 11, 23, 18, 23, 19, 13, 11, 10, 8, 8, 22, 4, 8, 21, 13, 9, 8, 6, 19, 6, 10, 10, 9, 9, 24, 22, 19, 15, 19, 6, 20, 6, 24, 19, 14, 17, 23, 9, 20, 20, 21, 18, 8, 8, 8, 10, 11, 21, 6, 23, 21, 20, 8, 8, 10, 19, 20, 21, 15, 15, 13, 18, 15, 20, 21, 18, 21, 19, 14, 20, 23, 13, 15, 15, 13, 19, 13, 8, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 13, 21, 6, 13, 19, 15, 17, 17, 13, 17, 15, 19, 6, 20, 13, 15, 14, 15, 21, 9, 23, 24, 18, 15, 15, 15, 19, 15, 15, 15, 17, 15, 13, 13, 15, 19, 14, 14, 14, 14, 14, 14, 20, 6, 11, 22, 21, 8, 9, 6, 17, 19, 6, 13, 19, 14, 19, 15, 13, 6, 11, 23, 9, 6, 14, 11, 15, 14, 15, 17, 19, 15, 14, 14, 15, 15, 14, 19, 19, 14, 15, 9, 15, 15, 6, 21, 20, 23, 23, 23, 23, 11, 19, 14, 19, 13, 9, 19, 19, 17, 23, 15, 15, 17, 14, 15, 15, 19, 13, 19, 22, 16, 25, 26, 27, 14, 15, 13, 15, 19, 13, 17, 14, 17, 14, 13, 11, 6, 9, 19, 15, 13, 6, 9, 19, 9, 19, 11, 20, 21, 19, 20, 24, 8, 10, 10, 11, 15, 13, 21, 8, 4, 23, 13, 17, 11, 15, 6, 8, 9, 24, 23, 6, 19, 10, 4, 11, 17, 17, 4, 8, 8, 9, 16, 24, 8, 17, 14, 23, 9, 6, 20, 16, 19, 9, 17, 23, 8, 23, 23, 23, 8, 8, 23, 9, 13, 6, 20, 23, 20, 4, 4, 8, 10, 8, 13, 20, 15, 11, 15, 19, 21, 6, 23, 11, 11, 11, 21, 15, 21, 23, 13, 19, 11, 23, 20, 11, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 4, 19, 13, 13, 20, 21, 13, 15, 15, 13, 21, 21, 15, 14, 19, 13, 14, 19, 15, 21, 13, 21, 21, 13, 23, 18, 21, 19, 19, 15, 15, 9, 23, 15, 15, 15, 15, 17, 17, 14, 14, 14, 19, 19, 17, 17, 20, 23, 23, 23, 23, 21, 23, 11, 20, 19, 21, 19, 18, 6, 8, 23, 23, 13, 15, 18, 17, 17, 15, 14, 13, 15, 14, 15, 6, 9, 11, 13, 19, 19, 13, 23, 20, 13, 20, 11, 13, 15, 19, 15, 14, 20, 23, 21, 14, 15, 15, 17, 17, 11, 15, 13, 15, 14, 14, 15, 15, 19, 6, 6, 19, 17, 15, 13, 29, 7, 14, 19, 13, 13, 18, 20, 20, 18, 9, 21, 15, 13, 23, 13, 20, 20, 19, 6, 6, 17, 20, 9, 8, 21, 23, 6, 6, 19, 20, 11, 11, 19, 9, 23, 24, 8, 8, 4, 19, 11, 9, 11, 15, 11, 11, 11, 13, 17, 11, 8, 23, 15, 21, 6, 20, 9, 9, 24, 16, 9, 8, 15, 18, 6, 9, 21, 23, 23, 9, 8, 20, 4, 9, 9, 8, 8, 8, 8, 22, 21, 21, 11, 13, 18, 8, 4, 9, 13, 13, 16, 6, 19, 21, 21, 20, 21, 13, 9, 8, 9, 21, 14, 15, 23, 6, 20, 14, 11, 6, 24, 16, 14, 4, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 13, 16, 24, 22, 6, 11, 23, 11, 13, 21, 20, 23, 18, 11, 13, 13, 13, 18, 20, 11, 18, 15, 18, 21, 18, 11, 23, 23, 21, 15, 15, 18, 18, 14, 15, 17, 15, 17, 19, 14, 15, 17, 17, 14, 14, 18, 20, 13, 23, 21, 9, 6, 11, 6, 20, 15, 15, 9, 11, 20, 11, 11, 21, 20, 11, 15, 17, 14, 14, 14, 19, 14, 13, 6, 19, 14, 14, 13, 9, 13, 19, 18, 13, 9, 20, 13, 6, 13, 6, 6, 4, 20, 15, 15, 13, 6, 14, 14, 14, 15, 14, 15, 14, 14, 15, 14, 14, 14, 19, 14, 14, 14, 18, 16, 16, 14, 15, 14, 19, 11, 9, 21, 23, 6, 18, 19, 21, 9, 9, 4, 9, 9, 6, 19, 15, 8, 8, 9, 6, 20, 23, 8, 8, 21, 14, 15, 9, 23, 23, 8, 8, 22, 9, 19, 19, 6, 11, 15, 23, 9, 19, 6, 15, 15, 20, 23, 23, 23, 9, 9, 24, 24, 11, 24, 23, 21, 13, 13, 15, 13, 6, 23, 23, 8, 8, 8, 6, 21, 23, 8, 8, 9, 24, 24, 23, 6, 21, 14, 15, 19, 23, 11, 13, 11, 9, 4, 19, 20, 23, 19, 19, 9, 6, 11, 11, 15, 15, 13, 8, 6, 15, 23, 18, 20, 23, 15, 15, 8, 0, 2, 2, 2, 2),
		(2, 1, 1, 1, 1, 0, 12, 7, 15, 15, 16, 24, 22, 24, 9, 8, 20, 15, 19, 21, 13, 17, 15, 13, 19, 6, 20, 15, 20, 18, 23, 19, 21, 23, 20, 19, 18, 21, 9, 9, 13, 15, 14, 15, 14, 14, 13, 6, 17, 17, 19, 17, 15, 15, 13, 17, 13, 23, 6, 9, 23, 20, 14, 13, 6, 9, 6, 18, 19, 19, 11, 13, 14, 19, 17, 11, 14, 17, 11, 15, 14, 14, 14, 21, 21, 21, 18, 15, 13, 21, 20, 13, 15, 20, 9, 21, 23, 19, 13, 4, 9, 11, 11, 15, 14, 14, 14, 14, 13, 11, 11, 13, 13, 17, 14, 14, 15, 15, 17, 18, 14, 15, 15, 15, 14, 14, 14, 19, 19, 23, 11, 23, 6, 6, 15, 11, 8, 9, 9, 23, 14, 9, 8, 24, 9, 6, 19, 4, 9, 6, 15, 23, 6, 15, 9, 8, 8, 10, 9, 19, 15, 18, 23, 9, 21, 15, 6, 9, 6, 14, 11, 21, 20, 6, 4, 23, 4, 24, 6, 4, 4, 19, 15, 23, 20, 15, 21, 23, 11, 23, 8, 4, 11, 15, 4, 8, 9, 6, 13, 19, 18, 19, 15, 15, 13, 11, 18, 23, 9, 20, 11, 9, 6, 18, 23, 23, 19, 20, 20, 6, 19, 14, 11, 9, 20, 21, 20, 13, 20, 9, 18, 14, 16, 7, 12, 0, 1, 1, 1, 1),
		(0, 1, 1, 1, 1, 2, 26, 26, 27, 28, 25, 16, 14, 16, 8, 24, 19, 19, 18, 15, 19, 14, 13, 13, 15, 23, 19, 21, 13, 11, 11, 13, 21, 13, 18, 15, 21, 6, 8, 9, 11, 15, 13, 15, 14, 14, 19, 17, 15, 15, 13, 13, 11, 17, 17, 14, 15, 19, 20, 20, 23, 15, 14, 13, 6, 23, 11, 11, 18, 15, 18, 20, 18, 9, 6, 19, 15, 15, 13, 15, 14, 13, 9, 20, 13, 21, 14, 15, 19, 11, 11, 20, 18, 18, 18, 9, 20, 21, 23, 20, 19, 15, 15, 17, 13, 17, 15, 17, 15, 24, 9, 19, 19, 13, 11, 17, 18, 22, 16, 7, 27, 28, 14, 17, 13, 20, 14, 15, 11, 20, 11, 9, 11, 9, 20, 19, 20, 21, 20, 14, 17, 11, 18, 16, 24, 11, 20, 9, 20, 15, 11, 20, 11, 19, 18, 20, 23, 9, 9, 11, 15, 21, 9, 9, 8, 13, 11, 9, 15, 5, 10, 4, 18, 9, 8, 6, 21, 9, 9, 4, 9, 19, 21, 19, 20, 13, 11, 20, 11, 11, 13, 17, 17, 15, 23, 23, 21, 17, 17, 17, 11, 9, 20, 11, 4, 9, 6, 18, 15, 23, 20, 6, 11, 19, 20, 18, 13, 11, 21, 20, 13, 6, 11, 13, 15, 19, 6, 24, 14, 16, 25, 28, 27, 26, 26, 2, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 28, 27, 26, 26, 26, 26, 27, 25, 16, 18, 19, 11, 20, 20, 19, 14, 11, 9, 14, 19, 19, 15, 21, 21, 19, 15, 19, 20, 20, 11, 6, 6, 14, 15, 19, 11, 19, 14, 13, 23, 11, 15, 14, 14, 17, 13, 19, 21, 15, 21, 19, 15, 15, 19, 13, 15, 15, 17, 6, 13, 13, 21, 23, 11, 13, 9, 22, 22, 13, 11, 6, 14, 14, 19, 11, 13, 23, 11, 13, 17, 15, 11, 11, 13, 21, 18, 21, 23, 19, 17, 17, 17, 17, 17, 19, 22, 16, 8, 9, 18, 8, 13, 15, 16, 18, 15, 21, 13, 9, 11, 16, 14, 14, 25, 26, 27, 18, 8, 6, 23, 11, 14, 14, 21, 6, 11, 13, 22, 24, 8, 22, 14, 14, 14, 11, 20, 21, 16, 11, 6, 18, 21, 13, 6, 4, 20, 11, 4, 11, 19, 19, 13, 9, 23, 13, 21, 19, 9, 4, 13, 21, 13, 21, 10, 10, 8, 19, 6, 10, 11, 23, 20, 13, 19, 19, 5, 13, 19, 6, 20, 20, 19, 6, 11, 19, 13, 13, 13, 13, 13, 13, 21, 24, 24, 9, 11, 23, 9, 9, 9, 8, 24, 16, 23, 13, 11, 11, 6, 19, 15, 23, 4, 9, 21, 20, 24, 24, 15, 15, 14, 15, 25, 27, 26, 26, 26, 26, 27, 28, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 5, 14, 14, 7, 25, 27, 26, 26, 27, 25, 14, 15, 16, 23, 19, 15, 14, 13, 14, 15, 19, 14, 15, 15, 19, 18, 20, 9, 23, 23, 9, 23, 14, 13, 9, 14, 14, 15, 19, 4, 13, 18, 13, 11, 14, 14, 15, 15, 20, 6, 6, 23, 13, 19, 15, 19, 15, 14, 15, 13, 11, 18, 6, 4, 4, 9, 19, 19, 4, 11, 13, 15, 15, 11, 23, 13, 15, 11, 15, 17, 15, 13, 13, 11, 23, 8, 4, 4, 6, 19, 13, 15, 18, 18, 20, 24, 9, 6, 11, 20, 23, 20, 15, 15, 13, 23, 21, 15, 21, 20, 9, 15, 14, 25, 26, 27, 16, 5, 11, 9, 6, 21, 23, 21, 15, 20, 13, 15, 11, 24, 13, 14, 15, 19, 6, 23, 9, 11, 13, 21, 15, 13, 9, 9, 22, 6, 13, 20, 9, 20, 11, 13, 23, 13, 6, 9, 15, 6, 20, 23, 19, 21, 8, 8, 9, 13, 4, 9, 21, 8, 9, 6, 21, 21, 15, 15, 15, 15, 11, 19, 13, 4, 13, 23, 9, 6, 19, 13, 21, 4, 4, 8, 9, 9, 24, 22, 8, 8, 9, 8, 24, 24, 10, 8, 23, 11, 17, 17, 14, 9, 4, 23, 18, 20, 23, 22, 18, 15, 14, 25, 27, 26, 26, 27, 28, 7, 14, 14, 5, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 4, 13, 15, 15, 14, 14, 5, 28, 26, 26, 26, 25, 14, 15, 17, 15, 15, 15, 14, 15, 17, 15, 19, 19, 21, 18, 20, 23, 13, 13, 13, 19, 11, 6, 19, 14, 8, 21, 19, 14, 15, 13, 6, 6, 13, 15, 14, 15, 21, 13, 23, 6, 9, 11, 18, 15, 17, 17, 14, 18, 19, 6, 23, 9, 9, 9, 17, 14, 17, 17, 19, 13, 14, 17, 11, 6, 19, 14, 20, 24, 16, 24, 9, 6, 23, 9, 6, 13, 13, 9, 22, 8, 10, 24, 15, 15, 13, 19, 15, 23, 13, 13, 11, 18, 15, 11, 20, 11, 14, 11, 18, 11, 15, 25, 26, 27, 14, 22, 4, 9, 13, 23, 10, 9, 11, 21, 15, 13, 6, 14, 19, 18, 14, 23, 11, 19, 6, 9, 6, 18, 18, 4, 4, 11, 8, 8, 9, 23, 8, 8, 18, 20, 20, 14, 21, 6, 11, 14, 13, 9, 19, 19, 9, 8, 24, 13, 10, 9, 13, 23, 8, 9, 15, 14, 18, 19, 6, 6, 18, 11, 11, 11, 13, 23, 6, 15, 13, 23, 23, 8, 8, 8, 9, 9, 24, 10, 8, 8, 10, 9, 21, 8, 10, 9, 13, 15, 11, 13, 14, 6, 8, 13, 11, 23, 23, 14, 14, 25, 26, 26, 26, 28, 10, 16, 16, 16, 15, 18, 4, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 18, 14, 15, 19, 21, 21, 15, 13, 25, 26, 26, 27, 29, 14, 19, 17, 15, 19, 15, 19, 13, 6, 11, 20, 15, 21, 11, 18, 18, 19, 23, 23, 21, 15, 20, 8, 23, 21, 15, 23, 11, 13, 17, 17, 11, 19, 9, 23, 15, 15, 21, 15, 19, 9, 13, 14, 15, 14, 21, 19, 19, 13, 20, 20, 19, 17, 14, 15, 15, 15, 17, 13, 15, 13, 11, 20, 19, 24, 8, 24, 24, 11, 19, 9, 9, 11, 15, 23, 8, 8, 24, 8, 8, 6, 13, 17, 14, 14, 19, 11, 11, 23, 18, 23, 9, 21, 21, 9, 20, 13, 11, 19, 17, 29, 5, 14, 20, 24, 13, 9, 6, 6, 9, 6, 13, 15, 14, 14, 13, 6, 21, 23, 20, 23, 9, 21, 19, 13, 13, 6, 21, 9, 4, 9, 9, 8, 9, 23, 8, 9, 18, 9, 6, 23, 20, 11, 18, 9, 8, 11, 14, 6, 8, 21, 13, 17, 13, 23, 18, 13, 15, 15, 6, 8, 9, 8, 8, 21, 21, 15, 20, 9, 21, 19, 13, 9, 8, 20, 20, 8, 8, 8, 9, 10, 10, 8, 8, 8, 22, 9, 8, 22, 9, 9, 17, 13, 15, 6, 21, 18, 6, 6, 16, 14, 29, 27, 26, 26, 25, 11, 16, 24, 8, 6, 19, 6, 24, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 22, 19, 14, 19, 11, 11, 23, 22, 15, 15, 28, 26, 26, 28, 15, 14, 17, 17, 19, 19, 18, 20, 20, 6, 13, 15, 15, 15, 17, 17, 6, 17, 15, 17, 13, 17, 19, 11, 23, 13, 20, 20, 23, 11, 19, 15, 19, 11, 11, 13, 15, 19, 8, 6, 15, 19, 15, 14, 15, 11, 11, 11, 13, 15, 15, 17, 14, 17, 11, 14, 14, 23, 20, 15, 13, 22, 9, 21, 6, 20, 9, 19, 23, 9, 19, 20, 9, 8, 8, 4, 6, 20, 20, 11, 13, 14, 15, 14, 13, 11, 23, 21, 23, 21, 20, 20, 13, 11, 19, 5, 23, 20, 18, 16, 14, 14, 20, 21, 23, 9, 13, 13, 23, 11, 21, 17, 14, 17, 19, 13, 15, 6, 9, 24, 23, 10, 24, 21, 13, 6, 15, 11, 8, 10, 10, 9, 8, 4, 8, 9, 11, 15, 9, 4, 11, 19, 13, 6, 11, 17, 13, 13, 11, 15, 21, 20, 11, 21, 20, 14, 19, 4, 4, 4, 23, 13, 18, 9, 6, 8, 9, 11, 17, 14, 6, 9, 6, 9, 13, 4, 9, 24, 8, 10, 8, 8, 8, 22, 13, 9, 11, 8, 10, 10, 24, 17, 15, 21, 20, 11, 11, 14, 14, 28, 26, 26, 28, 22, 14, 22, 4, 6, 11, 11, 6, 9, 11, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 13, 20, 23, 14, 18, 19, 13, 13, 21, 20, 16, 7, 27, 26, 27, 4, 16, 21, 18, 22, 8, 9, 11, 6, 13, 17, 15, 14, 15, 13, 13, 14, 13, 13, 14, 14, 17, 6, 23, 21, 14, 13, 23, 23, 15, 18, 18, 14, 13, 11, 15, 15, 15, 13, 17, 9, 11, 19, 15, 14, 6, 17, 14, 13, 11, 15, 14, 18, 13, 20, 13, 13, 21, 11, 15, 23, 9, 20, 14, 13, 13, 20, 11, 19, 11, 9, 8, 23, 23, 23, 11, 21, 15, 11, 11, 13, 11, 14, 6, 4, 23, 15, 15, 15, 21, 6, 6, 19, 11, 15, 20, 8, 22, 14, 15, 14, 15, 13, 9, 20, 19, 20, 6, 13, 18, 19, 13, 11, 11, 15, 19, 6, 9, 8, 24, 22, 8, 8, 6, 24, 13, 4, 9, 8, 10, 9, 24, 8, 9, 6, 23, 18, 23, 9, 21, 11, 21, 15, 19, 13, 11, 13, 17, 19, 20, 23, 20, 23, 18, 15, 16, 6, 8, 4, 8, 13, 15, 8, 4, 13, 19, 10, 10, 20, 13, 11, 20, 13, 21, 9, 24, 8, 8, 8, 10, 10, 9, 16, 22, 24, 4, 8, 8, 8, 23, 19, 14, 14, 16, 13, 15, 5, 27, 26, 27, 7, 16, 20, 21, 20, 21, 11, 20, 11, 11, 21, 11, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 16, 20, 11, 21, 15, 20, 13, 20, 15, 24, 18, 15, 15, 25, 26, 26, 25, 14, 14, 6, 5, 8, 9, 13, 15, 17, 13, 13, 17, 18, 15, 6, 4, 9, 15, 9, 9, 9, 11, 18, 18, 15, 13, 15, 11, 9, 9, 13, 21, 14, 14, 18, 15, 19, 15, 13, 17, 13, 6, 15, 14, 14, 14, 15, 13, 6, 13, 19, 13, 11, 11, 13, 18, 19, 19, 17, 19, 9, 13, 15, 20, 23, 21, 6, 9, 21, 21, 19, 19, 19, 11, 11, 13, 11, 9, 4, 20, 14, 17, 6, 21, 20, 21, 15, 14, 14, 14, 9, 11, 19, 15, 16, 29, 27, 28, 15, 15, 14, 15, 13, 6, 6, 4, 21, 18, 6, 9, 18, 11, 15, 15, 15, 8, 8, 9, 9, 8, 24, 5, 10, 8, 24, 8, 9, 8, 10, 9, 6, 19, 16, 13, 15, 21, 15, 11, 8, 8, 19, 14, 11, 13, 14, 14, 6, 8, 8, 6, 13, 15, 6, 9, 11, 8, 4, 13, 15, 13, 21, 11, 6, 13, 10, 23, 9, 23, 8, 4, 23, 19, 18, 16, 9, 10, 4, 8, 11, 13, 9, 8, 8, 8, 8, 8, 20, 11, 15, 14, 22, 24, 14, 25, 26, 26, 25, 15, 16, 22, 8, 20, 11, 15, 19, 11, 9, 21, 20, 13, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 16, 11, 11, 23, 20, 13, 23, 18, 15, 17, 14, 11, 22, 14, 29, 26, 26, 28, 14, 15, 11, 20, 20, 13, 17, 13, 19, 19, 13, 20, 20, 23, 23, 24, 16, 8, 8, 15, 15, 11, 9, 9, 16, 8, 4, 9, 9, 9, 14, 15, 8, 6, 21, 19, 15, 17, 19, 19, 17, 14, 15, 17, 13, 19, 15, 11, 20, 15, 11, 20, 19, 15, 18, 14, 15, 14, 19, 13, 18, 14, 18, 19, 19, 13, 13, 13, 11, 13, 13, 11, 9, 23, 23, 19, 23, 23, 20, 13, 15, 15, 15, 9, 11, 15, 14, 14, 11, 15, 18, 22, 6, 14, 25, 26, 27, 14, 16, 15, 18, 18, 11, 6, 19, 20, 9, 20, 24, 24, 24, 14, 17, 6, 21, 15, 8, 10, 9, 16, 10, 10, 8, 8, 8, 24, 22, 22, 11, 16, 6, 6, 18, 14, 23, 23, 9, 9, 11, 14, 15, 17, 15, 14, 15, 4, 9, 23, 11, 13, 9, 4, 4, 9, 13, 20, 19, 19, 19, 19, 24, 4, 19, 24, 23, 8, 8, 9, 4, 9, 11, 19, 8, 24, 16, 21, 16, 22, 6, 6, 8, 8, 8, 8, 9, 15, 17, 15, 15, 5, 22, 28, 26, 26, 29, 16, 22, 24, 11, 6, 13, 15, 11, 9, 20, 18, 11, 6, 11, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 22, 23, 6, 11, 23, 18, 13, 13, 17, 17, 17, 17, 19, 21, 16, 17, 27, 26, 28, 14, 16, 11, 13, 11, 24, 11, 19, 15, 15, 21, 9, 9, 11, 13, 6, 13, 19, 11, 9, 4, 8, 9, 20, 9, 4, 6, 20, 6, 19, 13, 9, 9, 23, 19, 13, 13, 17, 14, 14, 17, 6, 13, 24, 8, 9, 13, 19, 15, 19, 15, 13, 13, 11, 11, 17, 15, 14, 14, 14, 17, 14, 15, 23, 13, 20, 13, 13, 11, 6, 11, 23, 13, 19, 11, 23, 15, 15, 15, 13, 14, 19, 17, 13, 14, 15, 15, 20, 19, 9, 11, 19, 16, 25, 26, 27, 15, 16, 6, 23, 13, 17, 15, 15, 6, 11, 8, 8, 11, 14, 6, 6, 18, 21, 9, 13, 23, 9, 22, 8, 10, 8, 24, 8, 8, 24, 19, 20, 20, 9, 23, 18, 13, 23, 8, 20, 20, 6, 15, 17, 13, 14, 14, 14, 15, 6, 6, 24, 24, 8, 8, 9, 9, 21, 14, 13, 16, 22, 24, 24, 9, 4, 15, 9, 8, 8, 24, 23, 8, 13, 19, 11, 23, 9, 9, 13, 13, 19, 11, 4, 4, 9, 23, 18, 18, 9, 18, 24, 16, 28, 26, 27, 11, 16, 20, 11, 6, 6, 13, 19, 15, 13, 20, 11, 19, 20, 11, 6, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 24, 23, 13, 19, 20, 23, 18, 14, 17, 13, 19, 15, 13, 7, 19, 18, 14, 27, 26, 28, 14, 21, 13, 4, 8, 18, 15, 9, 15, 13, 11, 13, 13, 4, 13, 15, 13, 4, 8, 9, 6, 23, 10, 24, 19, 6, 4, 13, 6, 10, 13, 9, 6, 17, 14, 13, 17, 15, 6, 17, 14, 19, 20, 6, 6, 11, 14, 14, 14, 11, 11, 17, 19, 13, 14, 15, 14, 14, 14, 17, 11, 21, 13, 6, 6, 9, 9, 6, 9, 4, 9, 15, 21, 23, 13, 14, 14, 19, 13, 15, 15, 19, 14, 14, 13, 19, 14, 6, 11, 17, 15, 14, 29, 26, 27, 14, 22, 6, 9, 13, 17, 14, 17, 4, 11, 24, 23, 15, 19, 4, 11, 20, 11, 6, 9, 21, 15, 11, 8, 9, 8, 24, 9, 8, 9, 9, 21, 14, 18, 9, 19, 21, 20, 20, 23, 23, 11, 6, 19, 19, 13, 11, 13, 15, 13, 9, 24, 10, 10, 4, 8, 19, 14, 19, 17, 23, 8, 10, 8, 22, 9, 14, 8, 8, 8, 9, 11, 20, 9, 15, 19, 8, 10, 6, 9, 9, 6, 6, 19, 19, 20, 6, 16, 9, 11, 22, 16, 28, 26, 27, 16, 5, 23, 13, 11, 20, 16, 20, 13, 18, 20, 21, 18, 11, 23, 13, 16, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 21, 23, 6, 9, 23, 23, 20, 14, 15, 13, 19, 13, 17, 16, 11, 17, 18, 14, 27, 26, 28, 15, 9, 24, 24, 15, 11, 13, 21, 11, 18, 19, 9, 4, 18, 8, 20, 21, 4, 4, 13, 9, 24, 8, 24, 11, 23, 13, 8, 6, 20, 19, 9, 19, 15, 15, 13, 13, 13, 9, 23, 13, 17, 14, 17, 13, 6, 15, 13, 13, 14, 11, 17, 15, 15, 13, 19, 13, 14, 17, 20, 13, 14, 13, 9, 9, 8, 8, 8, 9, 6, 15, 23, 13, 18, 13, 19, 15, 13, 13, 17, 17, 14, 17, 13, 15, 14, 13, 15, 17, 17, 5, 5, 7, 17, 14, 14, 19, 15, 15, 15, 15, 19, 6, 21, 19, 21, 14, 17, 11, 13, 23, 4, 23, 6, 4, 8, 19, 23, 9, 6, 20, 9, 8, 10, 4, 13, 15, 18, 13, 17, 11, 15, 20, 9, 23, 19, 13, 20, 15, 20, 13, 6, 8, 23, 15, 9, 4, 4, 9, 19, 18, 9, 9, 11, 20, 8, 8, 8, 9, 13, 18, 24, 8, 8, 8, 11, 21, 9, 9, 20, 9, 20, 13, 9, 9, 6, 11, 23, 23, 20, 19, 16, 22, 11, 14, 28, 26, 27, 22, 23, 20, 6, 24, 18, 15, 23, 20, 13, 18, 11, 13, 19, 20, 19, 19, 13, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 24, 23, 13, 23, 9, 23, 18, 15, 15, 15, 11, 13, 19, 23, 17, 15, 23, 24, 14, 27, 26, 25, 22, 9, 16, 15, 15, 23, 6, 11, 9, 9, 21, 18, 23, 4, 8, 21, 9, 13, 18, 6, 8, 4, 4, 16, 15, 19, 20, 23, 9, 13, 15, 15, 11, 13, 11, 21, 24, 9, 22, 13, 11, 6, 17, 15, 19, 17, 19, 15, 15, 19, 15, 21, 8, 21, 19, 14, 14, 15, 15, 13, 23, 15, 6, 8, 9, 8, 8, 23, 15, 21, 6, 20, 23, 21, 19, 14, 11, 11, 15, 14, 15, 15, 14, 15, 15, 15, 17, 13, 20, 6, 20, 18, 15, 14, 11, 15, 14, 15, 23, 11, 17, 19, 16, 24, 20, 15, 14, 17, 23, 23, 8, 8, 9, 11, 9, 4, 13, 15, 17, 13, 8, 4, 22, 16, 13, 11, 18, 14, 15, 11, 13, 23, 8, 20, 19, 13, 8, 18, 18, 20, 8, 23, 20, 13, 11, 11, 16, 19, 20, 9, 4, 6, 6, 20, 22, 10, 8, 9, 11, 11, 22, 8, 22, 16, 9, 4, 6, 8, 21, 9, 13, 9, 19, 15, 13, 20, 9, 9, 9, 6, 6, 11, 14, 25, 26, 27, 16, 8, 10, 17, 5, 20, 6, 13, 20, 23, 11, 13, 13, 19, 21, 20, 11, 13, 16, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 23, 23, 13, 13, 11, 21, 18, 20, 18, 15, 13, 11, 17, 20, 19, 11, 11, 22, 18, 16, 27, 26, 29, 14, 17, 14, 23, 8, 17, 9, 6, 18, 11, 9, 20, 9, 4, 23, 13, 13, 6, 8, 24, 9, 6, 13, 18, 11, 8, 6, 11, 20, 18, 15, 23, 20, 15, 19, 13, 20, 23, 23, 20, 11, 18, 19, 17, 15, 14, 14, 15, 11, 11, 15, 13, 15, 19, 13, 13, 13, 19, 13, 21, 19, 20, 8, 9, 11, 20, 15, 15, 23, 23, 21, 23, 13, 15, 15, 15, 13, 14, 14, 16, 19, 15, 17, 14, 14, 14, 16, 16, 13, 6, 4, 11, 14, 14, 14, 14, 14, 15, 6, 17, 15, 22, 20, 14, 19, 20, 9, 11, 13, 9, 8, 10, 8, 22, 22, 9, 9, 20, 15, 18, 6, 6, 18, 21, 11, 17, 17, 6, 15, 13, 19, 10, 16, 24, 8, 23, 19, 13, 11, 23, 23, 20, 23, 11, 15, 19, 11, 11, 10, 4, 6, 11, 9, 23, 20, 8, 23, 23, 13, 14, 16, 22, 8, 8, 8, 20, 6, 6, 18, 13, 11, 16, 11, 9, 11, 21, 20, 13, 13, 9, 21, 7, 26, 26, 5, 16, 5, 6, 6, 13, 9, 8, 9, 13, 13, 11, 13, 15, 13, 11, 11, 8, 9, 13, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 4, 16, 13, 11, 11, 13, 15, 23, 13, 23, 23, 18, 13, 17, 13, 11, 23, 6, 5, 15, 16, 7, 26, 26, 16, 16, 15, 9, 21, 11, 9, 18, 11, 4, 10, 9, 23, 20, 11, 11, 6, 9, 11, 16, 24, 24, 4, 8, 9, 9, 20, 13, 13, 6, 18, 15, 21, 21, 17, 19, 6, 23, 23, 13, 15, 21, 11, 13, 14, 14, 15, 21, 18, 11, 13, 14, 14, 15, 6, 19, 6, 13, 23, 13, 18, 15, 13, 11, 13, 15, 19, 18, 20, 21, 21, 11, 19, 19, 11, 17, 15, 14, 19, 19, 22, 21, 14, 15, 7, 28, 27, 27, 26, 26, 26, 26, 27, 27, 27, 28, 25, 18, 14, 18, 15, 15, 15, 13, 13, 22, 8, 4, 23, 23, 6, 9, 24, 22, 11, 20, 23, 11, 18, 14, 15, 21, 21, 9, 6, 13, 13, 6, 13, 17, 15, 19, 11, 4, 24, 21, 19, 15, 11, 13, 19, 21, 21, 15, 20, 23, 11, 24, 4, 4, 6, 21, 9, 8, 13, 13, 13, 20, 13, 11, 15, 24, 10, 8, 8, 8, 13, 15, 15, 9, 9, 9, 4, 9, 9, 9, 11, 20, 11, 23, 16, 26, 26, 7, 16, 13, 6, 13, 13, 18, 6, 9, 6, 23, 13, 19, 14, 17, 11, 13, 21, 9, 6, 11, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 13, 13, 19, 11, 21, 21, 20, 21, 4, 8, 21, 15, 15, 11, 23, 13, 6, 6, 19, 24, 16, 29, 26, 27, 15, 16, 21, 20, 13, 19, 9, 4, 4, 4, 23, 9, 4, 20, 15, 15, 8, 8, 4, 11, 22, 4, 6, 9, 13, 8, 11, 20, 20, 15, 15, 18, 19, 11, 17, 11, 20, 23, 15, 15, 23, 19, 15, 15, 19, 17, 11, 18, 19, 19, 15, 6, 11, 19, 19, 13, 9, 13, 11, 11, 18, 19, 17, 15, 14, 15, 18, 19, 19, 11, 20, 15, 20, 11, 19, 14, 15, 11, 16, 17, 7, 28, 27, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 27, 29, 16, 14, 14, 17, 13, 18, 21, 23, 20, 11, 11, 17, 14, 15, 17, 19, 21, 15, 14, 15, 15, 14, 21, 9, 13, 14, 19, 13, 11, 22, 15, 14, 13, 21, 18, 20, 13, 14, 14, 14, 17, 15, 15, 23, 8, 23, 23, 4, 9, 22, 19, 20, 6, 9, 23, 15, 19, 8, 4, 13, 15, 22, 10, 8, 8, 9, 19, 15, 9, 4, 9, 8, 4, 9, 9, 11, 21, 4, 24, 14, 27, 26, 25, 16, 24, 13, 19, 20, 20, 19, 13, 13, 19, 21, 21, 11, 15, 19, 13, 11, 21, 20, 21, 19, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 16, 13, 23, 18, 15, 23, 19, 6, 6, 23, 23, 15, 13, 19, 13, 9, 9, 8, 24, 5, 17, 14, 28, 26, 25, 14, 4, 23, 15, 19, 9, 6, 11, 6, 20, 6, 6, 20, 9, 18, 9, 4, 4, 11, 11, 19, 13, 11, 11, 19, 19, 15, 15, 19, 6, 15, 19, 17, 15, 19, 18, 15, 15, 21, 19, 13, 13, 17, 17, 19, 20, 11, 15, 14, 15, 13, 11, 15, 21, 15, 13, 19, 14, 19, 13, 17, 14, 14, 17, 17, 15, 15, 21, 21, 15, 15, 15, 14, 19, 14, 15, 14, 7, 28, 26, 26, 26, 26, 26, 26, 27, 27, 28, 28, 28, 27, 27, 26, 26, 26, 26, 26, 26, 27, 29, 14, 14, 19, 15, 18, 19, 11, 23, 13, 17, 19, 13, 13, 21, 21, 13, 20, 20, 4, 6, 19, 18, 11, 17, 11, 8, 10, 22, 19, 17, 17, 13, 18, 9, 6, 17, 14, 13, 17, 17, 11, 9, 20, 23, 24, 24, 8, 24, 15, 13, 6, 6, 6, 20, 13, 9, 4, 13, 9, 22, 24, 8, 9, 24, 9, 4, 20, 4, 11, 9, 9, 24, 22, 15, 11, 19, 14, 25, 26, 27, 16, 11, 11, 13, 13, 20, 20, 11, 13, 20, 13, 21, 11, 19, 15, 15, 17, 11, 11, 21, 21, 16, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 24, 20, 23, 13, 18, 15, 21, 23, 11, 9, 23, 15, 15, 23, 20, 9, 4, 8, 20, 19, 6, 19, 16, 26, 26, 15, 16, 17, 11, 13, 15, 14, 15, 15, 19, 11, 13, 23, 9, 13, 19, 6, 17, 17, 17, 14, 19, 15, 21, 14, 15, 13, 13, 19, 19, 19, 15, 13, 19, 15, 15, 15, 17, 13, 17, 13, 11, 13, 18, 20, 9, 18, 13, 4, 23, 18, 9, 18, 21, 20, 14, 14, 14, 18, 13, 9, 11, 15, 17, 11, 11, 6, 20, 20, 15, 13, 21, 17, 17, 14, 15, 28, 26, 26, 26, 26, 27, 28, 29, 14, 16, 15, 14, 14, 16, 14, 15, 19, 29, 28, 27, 26, 26, 26, 26, 28, 17, 15, 17, 6, 19, 14, 14, 19, 13, 20, 6, 20, 19, 20, 23, 20, 19, 13, 9, 11, 15, 19, 15, 13, 8, 23, 20, 15, 15, 13, 19, 17, 17, 14, 15, 15, 14, 19, 13, 13, 20, 21, 20, 9, 24, 24, 6, 17, 19, 20, 8, 20, 20, 9, 23, 13, 6, 13, 23, 21, 9, 4, 23, 8, 8, 19, 20, 9, 24, 24, 11, 19, 13, 17, 15, 24, 26, 26, 5, 9, 6, 6, 20, 13, 15, 20, 20, 21, 24, 8, 24, 21, 15, 18, 15, 13, 15, 13, 9, 6, 11, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 24, 23, 21, 19, 11, 21, 14, 19, 23, 11, 15, 15, 6, 20, 9, 13, 6, 19, 15, 11, 11, 15, 18, 25, 26, 28, 14, 6, 15, 18, 15, 19, 19, 19, 19, 19, 11, 9, 11, 9, 23, 15, 15, 17, 15, 21, 20, 23, 13, 19, 13, 13, 13, 6, 9, 13, 21, 11, 11, 17, 14, 19, 11, 9, 19, 6, 9, 9, 6, 8, 11, 21, 9, 4, 9, 13, 23, 15, 15, 6, 20, 21, 20, 18, 13, 21, 11, 9, 15, 15, 18, 11, 23, 13, 21, 21, 13, 22, 14, 7, 27, 26, 26, 26, 27, 25, 14, 14, 16, 15, 14, 18, 19, 17, 19, 19, 6, 14, 20, 16, 18, 29, 27, 26, 26, 26, 26, 29, 14, 19, 6, 13, 13, 15, 18, 19, 11, 6, 8, 4, 4, 6, 21, 15, 20, 9, 8, 19, 19, 20, 13, 23, 20, 6, 11, 23, 15, 15, 5, 14, 14, 19, 15, 11, 13, 13, 15, 23, 23, 9, 24, 22, 19, 15, 20, 20, 21, 14, 20, 21, 21, 14, 19, 19, 20, 13, 17, 21, 23, 9, 11, 13, 14, 11, 24, 6, 17, 17, 15, 15, 16, 28, 26, 25, 21, 6, 9, 9, 9, 11, 18, 21, 21, 21, 11, 23, 21, 15, 13, 11, 18, 11, 18, 18, 20, 6, 19, 4, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 22, 21, 21, 18, 19, 19, 19, 21, 20, 13, 13, 23, 9, 11, 23, 9, 15, 19, 6, 19, 20, 13, 6, 14, 27, 26, 7, 14, 21, 11, 20, 21, 21, 11, 18, 14, 19, 6, 20, 9, 21, 14, 21, 23, 21, 9, 9, 21, 13, 9, 11, 16, 16, 9, 8, 24, 24, 6, 15, 17, 6, 21, 20, 18, 13, 11, 9, 6, 20, 20, 15, 9, 11, 9, 23, 4, 13, 19, 18, 23, 6, 21, 9, 23, 15, 14, 11, 20, 13, 14, 13, 20, 21, 13, 15, 19, 9, 15, 29, 26, 26, 26, 26, 25, 14, 16, 16, 6, 20, 17, 14, 14, 29, 27, 28, 18, 16, 17, 5, 5, 15, 14, 14, 29, 27, 26, 26, 26, 25, 14, 17, 13, 13, 13, 14, 15, 21, 21, 11, 9, 8, 6, 4, 19, 19, 21, 9, 13, 13, 19, 21, 20, 11, 4, 6, 15, 6, 9, 17, 14, 13, 9, 18, 23, 4, 6, 6, 8, 11, 20, 8, 4, 11, 15, 6, 8, 23, 21, 19, 18, 23, 23, 11, 21, 9, 9, 15, 19, 9, 23, 23, 11, 15, 13, 8, 13, 15, 15, 15, 18, 6, 26, 27, 15, 18, 23, 13, 18, 18, 18, 21, 18, 13, 20, 14, 15, 14, 19, 11, 13, 18, 21, 20, 19, 14, 14, 14, 4, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 24, 18, 15, 15, 18, 20, 11, 11, 15, 15, 23, 23, 9, 8, 15, 13, 23, 13, 19, 15, 9, 21, 17, 14, 29, 26, 28, 14, 23, 6, 24, 22, 22, 23, 15, 23, 9, 21, 15, 18, 15, 21, 9, 9, 23, 9, 15, 21, 11, 8, 10, 9, 18, 22, 24, 9, 22, 19, 15, 19, 6, 8, 20, 20, 8, 20, 13, 6, 15, 15, 13, 23, 11, 11, 21, 11, 13, 18, 19, 21, 23, 6, 13, 23, 14, 15, 13, 15, 21, 21, 20, 9, 13, 15, 17, 24, 15, 29, 26, 26, 26, 27, 6, 16, 18, 19, 7, 6, 11, 22, 19, 14, 25, 26, 26, 15, 16, 11, 18, 5, 6, 14, 14, 16, 15, 28, 26, 26, 26, 28, 14, 15, 13, 17, 20, 6, 13, 20, 13, 13, 6, 8, 8, 21, 8, 9, 21, 14, 11, 19, 13, 23, 20, 11, 20, 14, 9, 11, 14, 20, 9, 4, 23, 18, 13, 11, 6, 20, 9, 9, 8, 9, 13, 13, 23, 9, 13, 6, 20, 23, 23, 8, 4, 18, 6, 13, 6, 21, 23, 24, 23, 20, 23, 18, 22, 16, 17, 17, 23, 16, 28, 26, 25, 24, 6, 22, 18, 23, 11, 6, 13, 15, 15, 18, 15, 13, 17, 17, 21, 13, 15, 11, 13, 18, 15, 21, 19, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 22, 19, 14, 17, 6, 19, 11, 20, 13, 9, 21, 23, 6, 9, 13, 15, 6, 6, 14, 15, 11, 15, 15, 15, 14, 27, 26, 22, 16, 6, 11, 11, 6, 20, 23, 9, 6, 19, 15, 18, 13, 4, 13, 19, 21, 20, 13, 11, 23, 23, 9, 9, 17, 13, 23, 20, 18, 13, 15, 14, 13, 11, 18, 18, 23, 23, 20, 11, 15, 20, 23, 11, 13, 19, 20, 13, 15, 15, 13, 14, 13, 13, 13, 14, 18, 17, 13, 6, 17, 15, 15, 13, 19, 14, 15, 15, 29, 26, 26, 26, 28, 14, 16, 23, 6, 19, 17, 13, 13, 16, 15, 14, 25, 26, 27, 14, 16, 13, 18, 21, 21, 19, 15, 17, 15, 14, 25, 26, 26, 26, 28, 14, 19, 11, 20, 23, 23, 20, 6, 6, 11, 11, 18, 13, 9, 4, 9, 15, 15, 19, 15, 19, 19, 13, 15, 14, 13, 19, 11, 23, 23, 20, 4, 13, 20, 19, 23, 9, 4, 9, 11, 9, 19, 11, 11, 15, 6, 4, 23, 24, 9, 22, 20, 23, 19, 15, 9, 24, 22, 9, 9, 8, 4, 15, 17, 6, 21, 6, 24, 5, 26, 27, 16, 9, 13, 17, 11, 6, 6, 23, 19, 14, 18, 13, 19, 18, 11, 6, 11, 17, 14, 15, 15, 19, 20, 19, 16, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 14, 19, 9, 21, 20, 13, 20, 6, 6, 4, 20, 18, 19, 13, 23, 20, 19, 15, 19, 14, 15, 15, 13, 11, 16, 25, 26, 28, 16, 6, 6, 9, 23, 19, 13, 15, 20, 23, 15, 20, 11, 20, 15, 14, 20, 11, 6, 9, 9, 23, 20, 17, 17, 13, 18, 19, 18, 15, 15, 13, 15, 14, 9, 6, 20, 9, 21, 15, 13, 19, 23, 6, 23, 21, 11, 11, 13, 21, 23, 19, 19, 19, 19, 14, 23, 13, 15, 11, 13, 19, 17, 14, 14, 21, 16, 7, 26, 26, 26, 28, 14, 19, 4, 6, 6, 19, 15, 19, 17, 13, 13, 14, 25, 26, 27, 14, 19, 6, 16, 19, 9, 18, 13, 14, 15, 23, 16, 25, 26, 26, 26, 25, 14, 18, 20, 23, 9, 6, 18, 13, 4, 9, 20, 23, 13, 11, 19, 19, 6, 13, 14, 19, 11, 13, 14, 19, 14, 11, 8, 8, 9, 6, 21, 13, 6, 8, 11, 18, 23, 4, 13, 15, 15, 19, 24, 11, 11, 22, 8, 6, 9, 4, 8, 20, 18, 11, 24, 8, 24, 11, 11, 4, 13, 19, 17, 15, 20, 23, 16, 28, 26, 25, 16, 9, 20, 6, 6, 11, 13, 21, 19, 19, 15, 13, 19, 15, 20, 20, 15, 15, 15, 15, 11, 11, 19, 14, 16, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 15, 22, 8, 8, 21, 19, 21, 23, 9, 11, 18, 20, 15, 15, 11, 20, 19, 14, 14, 14, 19, 17, 6, 23, 8, 16, 26, 27, 16, 24, 6, 20, 18, 21, 13, 11, 6, 18, 14, 6, 13, 21, 18, 18, 11, 13, 11, 23, 9, 9, 20, 15, 14, 19, 15, 14, 15, 9, 9, 22, 22, 15, 19, 9, 6, 21, 18, 18, 9, 13, 23, 6, 9, 13, 11, 9, 23, 20, 22, 13, 19, 20, 15, 23, 11, 4, 8, 14, 19, 6, 19, 14, 14, 14, 15, 27, 26, 26, 28, 15, 16, 5, 6, 20, 20, 15, 15, 15, 13, 13, 19, 16, 14, 7, 11, 14, 11, 6, 21, 21, 13, 14, 11, 14, 15, 5, 24, 16, 25, 26, 26, 26, 29, 14, 15, 11, 11, 6, 13, 18, 19, 19, 9, 9, 19, 21, 15, 13, 20, 13, 19, 13, 15, 14, 17, 15, 19, 11, 23, 20, 13, 23, 11, 11, 20, 9, 9, 9, 20, 19, 20, 21, 20, 4, 8, 10, 8, 9, 9, 9, 4, 8, 8, 23, 13, 13, 17, 9, 13, 11, 17, 19, 13, 13, 15, 15, 6, 24, 16, 27, 26, 16, 10, 23, 11, 9, 11, 11, 20, 13, 20, 11, 15, 21, 21, 14, 19, 13, 19, 11, 11, 19, 6, 6, 18, 15, 16, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 6, 8, 22, 24, 9, 18, 15, 19, 13, 13, 21, 19, 21, 11, 21, 18, 14, 14, 13, 15, 9, 6, 17, 11, 24, 15, 28, 26, 7, 16, 23, 15, 21, 20, 13, 13, 11, 15, 21, 13, 13, 11, 21, 6, 19, 20, 11, 13, 13, 21, 21, 13, 17, 19, 21, 15, 19, 4, 8, 16, 8, 9, 13, 11, 13, 15, 18, 21, 23, 11, 6, 13, 9, 9, 11, 9, 23, 11, 24, 4, 24, 18, 13, 20, 11, 4, 23, 20, 18, 19, 15, 11, 11, 14, 28, 26, 26, 27, 14, 15, 19, 19, 18, 21, 19, 15, 19, 6, 13, 13, 13, 23, 19, 15, 15, 15, 17, 15, 23, 14, 14, 13, 6, 11, 15, 11, 9, 24, 18, 28, 26, 26, 27, 16, 15, 15, 17, 13, 23, 11, 15, 18, 6, 6, 18, 13, 15, 21, 19, 19, 14, 14, 15, 15, 13, 13, 17, 15, 13, 20, 6, 9, 10, 4, 11, 11, 9, 23, 19, 20, 6, 15, 20, 4, 24, 24, 10, 10, 16, 24, 4, 9, 23, 23, 11, 11, 15, 17, 6, 15, 15, 17, 6, 15, 13, 11, 21, 22, 29, 26, 28, 16, 8, 21, 6, 6, 13, 23, 9, 8, 23, 11, 19, 21, 19, 13, 19, 13, 13, 11, 19, 13, 23, 20, 18, 20, 15, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 9, 8, 9, 23, 9, 18, 13, 14, 13, 6, 18, 21, 6, 23, 21, 14, 15, 23, 19, 21, 9, 4, 13, 18, 11, 20, 29, 26, 28, 14, 19, 15, 13, 20, 13, 23, 20, 17, 11, 13, 9, 11, 13, 13, 18, 11, 23, 11, 20, 11, 8, 11, 19, 9, 11, 22, 22, 13, 6, 13, 9, 4, 6, 18, 19, 19, 20, 20, 21, 21, 11, 20, 8, 13, 15, 6, 6, 9, 9, 10, 11, 15, 9, 20, 20, 21, 23, 4, 14, 14, 19, 20, 19, 11, 26, 26, 26, 17, 21, 6, 15, 15, 15, 21, 15, 21, 18, 19, 13, 17, 22, 11, 16, 14, 15, 16, 17, 14, 14, 14, 15, 9, 22, 24, 21, 19, 6, 6, 24, 15, 27, 26, 26, 25, 15, 15, 17, 20, 22, 21, 22, 22, 14, 14, 13, 21, 13, 6, 23, 11, 11, 18, 15, 15, 15, 6, 13, 18, 20, 23, 9, 20, 8, 10, 9, 14, 13, 11, 9, 8, 4, 19, 19, 23, 20, 8, 23, 13, 20, 21, 23, 23, 16, 4, 9, 9, 9, 19, 14, 14, 19, 13, 14, 21, 13, 6, 15, 14, 28, 26, 4, 16, 13, 21, 11, 19, 21, 23, 6, 20, 21, 15, 18, 14, 19, 20, 15, 15, 17, 15, 15, 19, 20, 21, 21, 20, 14, 4, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 11, 8, 4, 8, 18, 21, 23, 21, 15, 15, 20, 9, 11, 23, 18, 15, 11, 19, 23, 21, 9, 8, 19, 15, 21, 24, 22, 26, 27, 14, 15, 13, 13, 23, 9, 13, 11, 21, 20, 20, 20, 14, 13, 11, 11, 19, 23, 13, 9, 4, 4, 18, 6, 4, 24, 9, 8, 16, 21, 8, 23, 9, 11, 18, 21, 13, 20, 19, 19, 11, 23, 23, 20, 19, 18, 11, 20, 9, 4, 9, 18, 20, 11, 9, 11, 14, 20, 11, 14, 15, 11, 24, 14, 28, 26, 26, 25, 18, 13, 13, 15, 19, 19, 19, 21, 9, 23, 13, 13, 17, 16, 14, 29, 27, 28, 14, 15, 14, 14, 14, 15, 4, 11, 23, 13, 14, 15, 17, 21, 18, 4, 26, 26, 27, 6, 5, 22, 13, 11, 21, 21, 21, 18, 20, 21, 13, 11, 23, 23, 23, 6, 20, 11, 15, 14, 14, 21, 23, 4, 13, 21, 20, 20, 19, 6, 11, 17, 19, 23, 21, 20, 19, 13, 14, 18, 13, 11, 11, 23, 8, 23, 23, 4, 4, 4, 9, 4, 13, 21, 19, 21, 20, 9, 9, 20, 9, 23, 14, 27, 26, 15, 21, 6, 11, 9, 20, 13, 11, 11, 13, 20, 11, 21, 15, 11, 11, 21, 21, 13, 15, 13, 13, 20, 21, 23, 20, 18, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 22, 4, 4, 8, 21, 21, 13, 11, 15, 14, 20, 11, 23, 19, 15, 13, 13, 9, 23, 21, 18, 11, 19, 21, 9, 16, 15, 27, 26, 7, 16, 20, 13, 19, 13, 18, 21, 20, 23, 9, 20, 20, 11, 11, 11, 19, 20, 8, 9, 6, 18, 13, 4, 9, 8, 8, 8, 6, 11, 21, 13, 13, 23, 9, 15, 13, 11, 21, 15, 18, 13, 9, 21, 19, 6, 9, 11, 9, 8, 18, 6, 23, 11, 20, 21, 23, 15, 15, 15, 6, 15, 16, 7, 26, 26, 27, 15, 23, 6, 11, 14, 14, 15, 15, 13, 23, 23, 13, 17, 19, 16, 15, 25, 26, 27, 14, 15, 13, 14, 14, 14, 15, 15, 15, 15, 14, 14, 11, 8, 10, 16, 28, 26, 26, 28, 8, 22, 19, 19, 19, 14, 14, 6, 4, 23, 15, 21, 8, 11, 13, 23, 15, 15, 6, 9, 6, 15, 15, 11, 11, 11, 15, 15, 18, 20, 14, 15, 13, 15, 20, 13, 21, 6, 13, 23, 15, 21, 9, 9, 4, 23, 9, 4, 4, 4, 16, 20, 19, 11, 13, 14, 21, 20, 21, 20, 20, 22, 7, 26, 27, 15, 13, 11, 19, 19, 18, 19, 20, 11, 11, 20, 21, 15, 21, 21, 13, 13, 21, 13, 13, 13, 19, 21, 21, 13, 21, 21, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 13, 11, 11, 17, 13, 11, 19, 18, 19, 15, 18, 11, 15, 15, 21, 20, 20, 23, 11, 13, 18, 13, 15, 21, 11, 15, 14, 25, 26, 25, 18, 13, 21, 9, 14, 21, 13, 23, 8, 8, 23, 21, 21, 13, 11, 9, 13, 8, 6, 18, 20, 23, 4, 8, 10, 8, 22, 9, 6, 19, 15, 11, 23, 21, 23, 19, 20, 20, 15, 14, 15, 9, 21, 13, 8, 6, 23, 4, 19, 15, 6, 4, 11, 20, 6, 23, 18, 14, 17, 6, 11, 14, 28, 26, 26, 25, 15, 18, 19, 14, 14, 13, 20, 15, 15, 18, 21, 15, 14, 17, 13, 14, 29, 26, 27, 14, 22, 7, 19, 19, 15, 14, 17, 17, 13, 17, 15, 19, 24, 23, 8, 5, 26, 26, 27, 16, 20, 11, 17, 14, 15, 11, 13, 11, 11, 15, 6, 13, 13, 9, 11, 14, 19, 9, 11, 6, 21, 15, 14, 17, 15, 11, 8, 6, 11, 23, 17, 11, 23, 23, 18, 19, 20, 6, 13, 11, 13, 13, 23, 11, 23, 8, 11, 23, 22, 11, 15, 19, 19, 11, 23, 18, 13, 11, 21, 18, 18, 25, 26, 25, 18, 11, 13, 18, 13, 20, 11, 23, 23, 23, 23, 21, 18, 21, 14, 20, 11, 19, 15, 11, 13, 17, 19, 21, 14, 21, 13, 4, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 13, 21, 21, 9, 6, 9, 15, 14, 11, 11, 19, 14, 15, 19, 11, 23, 23, 23, 20, 11, 6, 17, 14, 15, 17, 22, 17, 7, 26, 28, 16, 4, 5, 18, 18, 13, 23, 9, 6, 11, 15, 20, 6, 23, 9, 9, 23, 15, 19, 24, 8, 21, 24, 10, 10, 8, 24, 8, 8, 11, 15, 19, 18, 19, 19, 15, 15, 20, 20, 15, 14, 11, 19, 20, 23, 20, 20, 23, 15, 20, 15, 20, 19, 13, 23, 19, 13, 14, 13, 22, 11, 14, 27, 26, 27, 14, 17, 14, 14, 14, 14, 13, 13, 13, 13, 15, 15, 15, 15, 13, 14, 14, 25, 26, 27, 17, 11, 13, 17, 17, 17, 14, 19, 9, 6, 20, 19, 21, 11, 9, 8, 14, 27, 26, 26, 7, 15, 17, 15, 14, 15, 11, 11, 13, 13, 19, 11, 15, 14, 11, 15, 15, 13, 11, 23, 21, 20, 13, 21, 8, 4, 8, 8, 9, 13, 6, 20, 21, 11, 11, 17, 15, 9, 24, 23, 9, 9, 23, 18, 19, 9, 8, 11, 17, 11, 11, 17, 13, 17, 5, 5, 13, 17, 13, 18, 14, 14, 28, 26, 7, 17, 24, 11, 13, 6, 9, 11, 23, 9, 9, 20, 19, 20, 21, 18, 20, 6, 20, 19, 23, 23, 21, 6, 13, 13, 20, 9, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 11, 20, 23, 9, 13, 21, 9, 9, 13, 15, 13, 14, 14, 13, 5, 9, 9, 23, 11, 19, 13, 15, 14, 14, 11, 24, 13, 15, 26, 27, 16, 11, 13, 19, 23, 13, 11, 6, 20, 15, 21, 4, 9, 8, 8, 9, 13, 15, 6, 9, 22, 13, 8, 9, 9, 9, 8, 9, 18, 13, 17, 14, 18, 9, 6, 9, 20, 15, 21, 9, 15, 14, 15, 19, 11, 18, 19, 14, 21, 21, 19, 19, 13, 15, 14, 18, 18, 15, 19, 13, 14, 7, 26, 26, 28, 15, 14, 15, 14, 15, 15, 6, 11, 19, 6, 13, 14, 14, 14, 14, 14, 16, 17, 19, 16, 15, 11, 15, 14, 14, 14, 19, 14, 18, 21, 21, 15, 14, 15, 19, 16, 14, 25, 26, 26, 25, 14, 14, 14, 14, 14, 14, 14, 15, 14, 14, 14, 17, 13, 14, 14, 11, 13, 19, 13, 15, 18, 21, 21, 15, 15, 13, 13, 15, 14, 14, 14, 14, 15, 14, 14, 14, 15, 18, 19, 14, 18, 15, 14, 19, 15, 14, 14, 14, 14, 14, 14, 14, 14, 15, 19, 15, 14, 15, 19, 14, 14, 27, 26, 14, 17, 16, 15, 18, 13, 13, 19, 19, 21, 11, 19, 21, 19, 15, 21, 15, 18, 18, 13, 13, 19, 15, 19, 14, 18, 18, 19, 4, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 11, 13, 6, 11, 18, 23, 8, 6, 17, 14, 19, 17, 15, 13, 9, 6, 20, 20, 23, 13, 15, 19, 23, 18, 16, 9, 11, 18, 27, 27, 15, 17, 18, 24, 13, 18, 15, 11, 6, 19, 6, 8, 23, 9, 9, 19, 11, 6, 21, 9, 17, 13, 5, 11, 20, 20, 20, 21, 20, 11, 17, 19, 21, 4, 8, 11, 9, 20, 18, 13, 17, 14, 14, 15, 11, 19, 14, 15, 21, 18, 15, 21, 13, 15, 15, 19, 11, 11, 13, 15, 14, 28, 26, 26, 25, 15, 6, 19, 15, 14, 6, 6, 17, 15, 17, 15, 14, 14, 15, 14, 11, 8, 16, 22, 24, 14, 19, 19, 18, 9, 23, 23, 20, 21, 19, 4, 6, 9, 13, 6, 8, 24, 7, 26, 26, 27, 14, 14, 14, 19, 17, 13, 17, 15, 15, 19, 19, 17, 13, 19, 15, 15, 15, 13, 21, 19, 13, 23, 23, 19, 13, 14, 15, 14, 21, 13, 21, 15, 15, 15, 14, 14, 19, 16, 23, 11, 6, 11, 20, 20, 21, 13, 11, 17, 13, 15, 14, 6, 11, 19, 23, 11, 20, 14, 14, 14, 14, 26, 27, 15, 11, 17, 21, 23, 23, 23, 6, 11, 6, 23, 20, 23, 18, 23, 6, 19, 19, 11, 20, 21, 21, 14, 18, 19, 9, 21, 18, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 19, 23, 6, 19, 23, 9, 20, 13, 17, 15, 15, 19, 17, 15, 19, 13, 8, 8, 23, 13, 15, 21, 20, 20, 21, 6, 13, 16, 27, 26, 11, 15, 21, 20, 21, 14, 21, 9, 11, 11, 9, 6, 11, 20, 15, 20, 9, 23, 19, 15, 15, 15, 17, 17, 9, 6, 15, 21, 23, 11, 17, 23, 19, 13, 13, 11, 20, 13, 13, 19, 14, 14, 15, 17, 17, 17, 15, 6, 13, 20, 23, 21, 20, 6, 19, 20, 23, 18, 18, 14, 16, 27, 26, 26, 15, 22, 13, 19, 13, 14, 15, 13, 15, 17, 14, 14, 11, 11, 6, 11, 17, 15, 14, 19, 16, 16, 14, 23, 9, 24, 22, 9, 19, 23, 13, 11, 11, 23, 19, 19, 17, 19, 14, 27, 26, 26, 15, 14, 15, 11, 11, 17, 13, 13, 14, 13, 17, 6, 14, 19, 11, 6, 17, 19, 21, 13, 11, 23, 23, 19, 23, 11, 18, 21, 23, 6, 9, 8, 15, 15, 14, 15, 13, 22, 23, 9, 23, 4, 20, 16, 6, 4, 6, 13, 17, 17, 20, 20, 6, 20, 23, 23, 24, 18, 14, 11, 13, 26, 27, 16, 17, 17, 20, 9, 8, 8, 9, 23, 9, 6, 23, 19, 21, 11, 23, 20, 21, 6, 21, 18, 8, 23, 11, 11, 9, 11, 19, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 4, 6, 20, 6, 6, 6, 21, 19, 11, 14, 18, 19, 15, 11, 23, 19, 11, 9, 11, 23, 13, 15, 18, 11, 11, 18, 19, 5, 16, 28, 26, 4, 18, 15, 20, 11, 19, 20, 20, 18, 6, 9, 9, 20, 19, 23, 9, 13, 13, 18, 14, 17, 21, 20, 23, 13, 15, 18, 21, 15, 19, 21, 18, 15, 21, 13, 11, 23, 23, 13, 13, 13, 17, 15, 17, 6, 14, 17, 6, 11, 23, 23, 15, 20, 6, 18, 6, 6, 14, 19, 11, 15, 27, 26, 27, 14, 15, 15, 15, 15, 14, 14, 15, 14, 14, 19, 11, 19, 19, 13, 22, 16, 11, 28, 27, 27, 7, 14, 17, 23, 21, 19, 11, 14, 15, 13, 14, 14, 15, 13, 19, 6, 13, 14, 28, 26, 26, 7, 15, 21, 20, 11, 20, 21, 23, 15, 19, 13, 11, 16, 24, 23, 4, 4, 11, 11, 8, 4, 9, 9, 18, 20, 19, 19, 19, 17, 6, 9, 6, 15, 19, 17, 6, 17, 13, 13, 13, 11, 6, 24, 8, 24, 20, 20, 11, 17, 17, 17, 15, 11, 11, 11, 8, 21, 19, 13, 16, 6, 26, 28, 16, 13, 15, 19, 8, 8, 8, 9, 23, 13, 11, 19, 19, 13, 20, 9, 21, 19, 20, 23, 23, 4, 23, 11, 13, 6, 20, 19, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 9, 19, 21, 21, 15, 21, 11, 15, 15, 11, 13, 9, 20, 9, 6, 20, 19, 20, 11, 19, 18, 19, 11, 23, 19, 15, 11, 18, 28, 26, 7, 16, 17, 15, 11, 15, 9, 20, 19, 20, 9, 21, 14, 13, 11, 18, 21, 19, 21, 19, 15, 13, 20, 20, 18, 11, 6, 9, 23, 23, 23, 20, 8, 4, 9, 23, 6, 6, 23, 22, 18, 15, 15, 19, 14, 15, 14, 15, 13, 19, 15, 19, 19, 19, 21, 13, 14, 15, 13, 11, 15, 26, 26, 27, 14, 16, 13, 6, 19, 14, 17, 14, 15, 6, 11, 13, 19, 13, 6, 16, 29, 26, 26, 26, 26, 26, 25, 14, 14, 15, 19, 11, 17, 14, 13, 6, 13, 19, 4, 13, 17, 19, 14, 25, 26, 26, 29, 15, 19, 18, 21, 23, 21, 14, 20, 17, 15, 13, 9, 9, 23, 20, 13, 11, 20, 21, 20, 6, 20, 20, 13, 11, 9, 11, 15, 19, 18, 18, 18, 14, 17, 13, 15, 17, 13, 15, 14, 15, 20, 23, 20, 15, 13, 15, 14, 15, 17, 15, 17, 13, 18, 19, 18, 20, 23, 18, 7, 26, 28, 14, 11, 13, 15, 20, 22, 22, 23, 20, 18, 19, 15, 20, 13, 15, 15, 19, 20, 23, 23, 20, 23, 20, 14, 14, 15, 18, 11, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 19, 11, 20, 14, 11, 9, 13, 13, 13, 23, 6, 11, 9, 13, 21, 19, 20, 18, 13, 11, 19, 18, 6, 23, 15, 19, 15, 18, 28, 26, 29, 22, 6, 22, 19, 18, 11, 13, 11, 18, 15, 15, 11, 23, 13, 23, 9, 11, 19, 11, 15, 8, 23, 20, 9, 9, 23, 20, 13, 23, 23, 13, 6, 13, 6, 13, 13, 9, 9, 22, 9, 20, 6, 17, 17, 19, 17, 19, 13, 13, 11, 23, 20, 18, 11, 14, 14, 15, 17, 15, 19, 26, 26, 28, 15, 19, 14, 15, 14, 19, 19, 14, 19, 13, 13, 11, 11, 13, 17, 14, 27, 26, 26, 26, 26, 26, 27, 14, 15, 20, 6, 9, 9, 19, 13, 6, 9, 22, 13, 13, 15, 17, 14, 25, 26, 26, 25, 16, 20, 21, 13, 20, 11, 13, 13, 4, 15, 19, 4, 10, 8, 9, 6, 19, 9, 4, 23, 19, 9, 4, 19, 8, 10, 10, 8, 24, 20, 23, 9, 15, 23, 9, 11, 15, 15, 20, 6, 18, 15, 13, 17, 17, 15, 17, 8, 8, 4, 9, 21, 15, 19, 11, 9, 24, 4, 22, 29, 26, 28, 18, 6, 9, 15, 21, 22, 22, 9, 23, 19, 6, 6, 19, 15, 13, 13, 20, 13, 19, 21, 21, 19, 15, 14, 13, 19, 20, 19, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 4, 22, 20, 13, 13, 11, 21, 20, 9, 21, 23, 13, 13, 11, 20, 21, 6, 20, 11, 15, 11, 18, 19, 6, 18, 15, 13, 13, 14, 28, 26, 25, 24, 5, 24, 15, 14, 20, 20, 6, 21, 15, 19, 23, 9, 9, 6, 13, 19, 13, 13, 19, 13, 20, 9, 6, 11, 19, 19, 11, 23, 23, 21, 11, 21, 18, 13, 21, 23, 6, 23, 9, 20, 17, 14, 11, 19, 11, 11, 15, 14, 21, 11, 21, 18, 15, 13, 14, 6, 6, 19, 7, 26, 26, 28, 16, 17, 14, 14, 19, 17, 17, 19, 19, 14, 15, 14, 15, 15, 14, 15, 26, 26, 26, 26, 26, 26, 26, 29, 14, 13, 13, 11, 24, 22, 16, 8, 24, 22, 16, 19, 14, 14, 16, 29, 26, 26, 25, 15, 19, 19, 19, 19, 13, 13, 13, 19, 13, 13, 22, 8, 8, 9, 4, 13, 9, 23, 20, 21, 20, 20, 13, 9, 10, 10, 8, 22, 20, 8, 23, 15, 23, 8, 9, 18, 20, 8, 8, 8, 15, 14, 14, 14, 17, 15, 8, 8, 23, 20, 9, 8, 19, 20, 9, 10, 10, 5, 25, 26, 25, 16, 10, 23, 11, 11, 9, 8, 8, 23, 13, 11, 20, 20, 23, 20, 11, 9, 9, 16, 11, 4, 11, 14, 15, 13, 23, 9, 24, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 19, 6, 9, 6, 11, 18, 4, 6, 13, 13, 15, 17, 11, 9, 23, 13, 17, 15, 6, 11, 15, 17, 19, 18, 21, 13, 5, 18, 25, 26, 29, 16, 11, 22, 13, 15, 13, 11, 6, 13, 13, 18, 20, 23, 6, 6, 17, 13, 13, 6, 17, 15, 6, 6, 6, 19, 17, 20, 11, 23, 23, 21, 11, 13, 15, 13, 6, 6, 6, 9, 4, 19, 17, 17, 18, 11, 11, 19, 15, 19, 15, 17, 13, 15, 11, 9, 15, 6, 13, 16, 13, 26, 26, 28, 14, 14, 17, 15, 14, 15, 15, 14, 17, 15, 14, 19, 19, 20, 6, 17, 26, 26, 26, 26, 26, 26, 26, 29, 15, 19, 13, 19, 20, 11, 15, 11, 9, 11, 23, 18, 14, 14, 11, 29, 26, 26, 25, 14, 17, 17, 13, 11, 11, 11, 13, 13, 18, 9, 9, 21, 4, 10, 4, 11, 4, 20, 20, 9, 19, 21, 6, 6, 10, 10, 22, 24, 8, 24, 9, 19, 19, 9, 19, 9, 23, 9, 23, 19, 15, 19, 11, 6, 13, 19, 13, 11, 20, 6, 18, 21, 23, 13, 19, 22, 8, 8, 25, 26, 25, 16, 10, 9, 11, 23, 11, 9, 21, 15, 15, 11, 24, 9, 8, 9, 8, 8, 24, 24, 11, 11, 15, 14, 19, 9, 8, 8, 6, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 20, 8, 6, 18, 13, 8, 9, 17, 15, 15, 17, 6, 6, 23, 23, 11, 13, 19, 11, 11, 14, 15, 15, 4, 24, 13, 11, 14, 25, 26, 29, 16, 9, 9, 13, 14, 17, 15, 13, 6, 9, 19, 21, 11, 9, 21, 20, 11, 9, 20, 21, 9, 21, 6, 19, 21, 23, 13, 6, 6, 11, 13, 11, 6, 20, 20, 9, 20, 13, 6, 9, 14, 14, 11, 15, 21, 21, 14, 17, 9, 6, 15, 14, 13, 4, 13, 14, 17, 6, 15, 11, 26, 26, 28, 14, 19, 14, 14, 14, 15, 17, 11, 11, 11, 13, 13, 20, 23, 20, 16, 27, 26, 26, 26, 26, 26, 27, 15, 9, 15, 19, 21, 6, 8, 13, 6, 4, 8, 13, 21, 23, 18, 14, 25, 26, 26, 25, 16, 20, 21, 20, 13, 19, 15, 21, 20, 15, 15, 11, 21, 13, 9, 9, 23, 19, 9, 4, 20, 21, 9, 6, 20, 10, 22, 24, 8, 24, 22, 11, 11, 19, 18, 23, 9, 13, 19, 11, 13, 11, 13, 8, 23, 11, 23, 19, 13, 23, 11, 13, 4, 4, 23, 9, 22, 21, 16, 29, 26, 28, 16, 13, 23, 21, 19, 18, 18, 19, 9, 9, 8, 8, 8, 8, 8, 8, 9, 6, 6, 21, 14, 14, 21, 13, 9, 8, 8, 6, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 4, 15, 11, 19, 21, 4, 4, 20, 14, 17, 23, 23, 6, 20, 23, 8, 8, 13, 19, 14, 17, 19, 14, 15, 11, 22, 19, 17, 16, 28, 26, 29, 24, 8, 24, 15, 14, 17, 13, 21, 23, 23, 23, 9, 23, 9, 24, 10, 8, 9, 20, 9, 8, 20, 9, 23, 8, 23, 23, 23, 6, 20, 23, 6, 9, 9, 20, 9, 20, 21, 17, 19, 14, 15, 9, 9, 19, 11, 11, 19, 4, 13, 14, 13, 13, 15, 14, 15, 14, 14, 14, 13, 26, 26, 28, 14, 22, 22, 19, 15, 15, 14, 11, 22, 24, 4, 13, 21, 11, 6, 24, 7, 27, 26, 26, 26, 27, 7, 14, 20, 11, 19, 13, 18, 13, 23, 13, 6, 9, 15, 23, 8, 9, 14, 25, 26, 26, 25, 22, 24, 24, 24, 8, 20, 20, 8, 23, 11, 19, 19, 4, 6, 13, 21, 21, 11, 9, 23, 13, 20, 21, 13, 19, 15, 13, 6, 11, 22, 6, 13, 14, 13, 15, 13, 13, 13, 13, 23, 23, 23, 8, 9, 23, 20, 20, 8, 23, 13, 21, 19, 11, 8, 9, 9, 9, 8, 16, 6, 26, 28, 18, 6, 14, 18, 15, 15, 19, 20, 8, 9, 8, 4, 9, 6, 9, 8, 9, 11, 17, 19, 14, 11, 11, 19, 11, 9, 24, 13, 4, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 14, 15, 15, 6, 6, 18, 13, 6, 13, 20, 23, 23, 23, 9, 8, 8, 9, 6, 15, 14, 14, 17, 15, 20, 9, 21, 5, 16, 27, 26, 13, 8, 9, 22, 13, 17, 15, 13, 6, 11, 9, 4, 10, 9, 18, 10, 10, 24, 24, 23, 9, 8, 8, 18, 8, 8, 8, 8, 6, 23, 11, 6, 11, 11, 23, 15, 13, 21, 23, 11, 14, 19, 20, 8, 23, 15, 13, 11, 17, 15, 14, 15, 17, 13, 14, 14, 15, 17, 15, 19, 19, 27, 26, 27, 14, 5, 9, 20, 19, 13, 15, 21, 22, 9, 24, 13, 21, 23, 9, 17, 15, 22, 25, 28, 28, 17, 17, 6, 23, 23, 21, 11, 15, 14, 21, 13, 4, 18, 18, 9, 9, 13, 15, 28, 26, 26, 8, 22, 8, 8, 8, 24, 18, 8, 23, 23, 9, 6, 20, 23, 4, 9, 15, 8, 6, 4, 11, 11, 9, 20, 6, 19, 17, 6, 9, 6, 11, 17, 14, 17, 16, 15, 23, 23, 13, 19, 21, 23, 8, 8, 20, 21, 20, 23, 8, 23, 15, 11, 6, 20, 13, 21, 15, 21, 11, 22, 6, 26, 28, 18, 6, 17, 19, 9, 21, 15, 23, 6, 20, 13, 6, 17, 11, 6, 13, 15, 17, 11, 13, 14, 9, 11, 17, 11, 11, 18, 19, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 19, 15, 15, 19, 15, 15, 6, 9, 9, 19, 23, 9, 6, 6, 20, 21, 20, 20, 4, 20, 15, 4, 23, 20, 9, 13, 6, 16, 27, 26, 11, 22, 19, 11, 19, 19, 24, 11, 4, 4, 20, 9, 4, 9, 24, 23, 9, 20, 8, 20, 9, 10, 8, 13, 9, 8, 9, 8, 8, 22, 16, 13, 21, 23, 23, 13, 11, 8, 9, 15, 14, 17, 19, 17, 14, 14, 14, 19, 15, 14, 19, 6, 6, 19, 13, 17, 14, 14, 14, 20, 15, 27, 26, 26, 16, 24, 13, 20, 23, 9, 21, 19, 13, 23, 18, 11, 6, 19, 17, 13, 16, 17, 16, 16, 13, 17, 23, 8, 8, 10, 8, 22, 20, 20, 18, 14, 14, 17, 15, 22, 19, 11, 16, 27, 26, 26, 8, 8, 8, 8, 10, 22, 23, 8, 9, 9, 8, 9, 9, 8, 6, 20, 23, 13, 19, 20, 11, 9, 9, 9, 20, 23, 20, 6, 11, 13, 15, 11, 13, 13, 24, 23, 13, 6, 11, 15, 13, 8, 9, 23, 20, 11, 9, 4, 6, 11, 6, 17, 11, 13, 23, 9, 17, 15, 23, 5, 11, 26, 27, 14, 6, 24, 6, 21, 19, 21, 23, 9, 6, 20, 11, 11, 11, 15, 14, 18, 21, 18, 14, 14, 11, 11, 15, 17, 14, 19, 19, 4, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 4, 16, 15, 19, 17, 13, 23, 23, 23, 8, 23, 18, 19, 19, 11, 20, 20, 8, 10, 10, 22, 22, 9, 3, 6, 18, 20, 9, 24, 26, 26, 16, 15, 13, 13, 15, 16, 8, 9, 4, 10, 23, 20, 11, 9, 10, 20, 15, 9, 9, 11, 9, 9, 23, 9, 19, 13, 23, 8, 8, 9, 4, 9, 20, 23, 6, 11, 14, 13, 15, 14, 19, 11, 15, 18, 21, 19, 20, 21, 15, 18, 13, 13, 15, 15, 17, 17, 15, 15, 14, 15, 18, 28, 26, 26, 25, 18, 5, 23, 23, 20, 6, 15, 15, 15, 6, 8, 6, 9, 20, 16, 6, 17, 5, 5, 16, 15, 23, 9, 10, 10, 21, 15, 23, 9, 9, 14, 14, 6, 13, 16, 17, 24, 13, 26, 26, 27, 16, 10, 8, 10, 5, 13, 8, 9, 9, 9, 8, 9, 9, 8, 15, 19, 8, 8, 19, 14, 4, 4, 9, 20, 13, 4, 20, 20, 19, 15, 17, 6, 17, 11, 8, 8, 19, 11, 20, 23, 13, 21, 20, 6, 23, 21, 20, 11, 13, 6, 8, 9, 20, 20, 23, 23, 11, 11, 11, 22, 14, 27, 26, 15, 6, 16, 23, 14, 21, 6, 19, 11, 11, 13, 19, 18, 15, 21, 6, 9, 11, 21, 20, 20, 13, 13, 15, 19, 6, 6, 20, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 4, 15, 19, 13, 6, 6, 9, 23, 11, 13, 20, 20, 19, 20, 6, 6, 23, 4, 10, 8, 22, 10, 11, 9, 20, 8, 8, 17, 9, 26, 27, 14, 6, 17, 19, 11, 11, 24, 6, 21, 4, 11, 24, 22, 9, 9, 6, 23, 11, 4, 20, 6, 19, 6, 9, 11, 20, 4, 10, 10, 24, 22, 19, 14, 18, 18, 18, 15, 19, 14, 11, 23, 8, 18, 13, 11, 21, 19, 15, 19, 11, 20, 14, 15, 13, 15, 15, 17, 13, 19, 17, 22, 29, 26, 26, 28, 14, 13, 15, 11, 20, 9, 20, 18, 9, 8, 23, 8, 10, 8, 16, 13, 22, 10, 25, 29, 14, 24, 4, 13, 19, 21, 19, 6, 9, 20, 13, 19, 17, 17, 19, 9, 20, 25, 26, 26, 28, 16, 6, 9, 13, 19, 11, 9, 11, 9, 9, 8, 9, 19, 16, 6, 21, 8, 10, 11, 20, 4, 4, 21, 18, 18, 9, 9, 11, 23, 13, 20, 23, 11, 8, 24, 24, 19, 15, 13, 23, 18, 15, 11, 23, 13, 23, 21, 11, 8, 23, 9, 9, 9, 21, 23, 11, 11, 17, 17, 13, 16, 27, 26, 19, 15, 20, 15, 15, 19, 13, 13, 19, 9, 21, 15, 20, 11, 9, 9, 6, 20, 13, 23, 23, 13, 11, 24, 22, 9, 6, 11, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 11, 14, 15, 13, 13, 6, 20, 9, 8, 10, 10, 9, 15, 15, 11, 8, 8, 8, 24, 24, 10, 4, 13, 19, 9, 8, 15, 4, 26, 28, 5, 9, 9, 19, 11, 11, 24, 9, 20, 20, 13, 20, 8, 19, 13, 4, 8, 20, 19, 23, 11, 9, 11, 9, 9, 18, 13, 22, 22, 21, 6, 11, 11, 9, 6, 23, 21, 14, 20, 8, 24, 21, 22, 19, 19, 19, 19, 14, 13, 19, 13, 17, 14, 17, 17, 15, 16, 13, 9, 11, 15, 15, 27, 26, 27, 16, 22, 15, 9, 23, 23, 8, 8, 23, 9, 22, 22, 10, 8, 13, 15, 16, 25, 26, 27, 14, 16, 17, 15, 17, 17, 6, 6, 11, 20, 4, 6, 19, 13, 17, 5, 16, 27, 26, 26, 4, 5, 5, 23, 11, 4, 17, 20, 13, 20, 11, 6, 6, 11, 9, 9, 9, 9, 20, 4, 9, 21, 21, 21, 9, 9, 23, 19, 21, 8, 9, 20, 23, 23, 20, 8, 22, 15, 15, 19, 19, 23, 11, 23, 13, 6, 20, 21, 6, 9, 9, 23, 24, 8, 23, 18, 20, 11, 17, 11, 5, 16, 28, 26, 10, 14, 14, 15, 19, 20, 19, 9, 13, 15, 19, 20, 9, 9, 6, 23, 11, 20, 11, 20, 20, 11, 6, 8, 22, 22, 22, 16, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 16, 17, 15, 15, 19, 13, 11, 10, 8, 8, 8, 20, 6, 15, 21, 9, 20, 22, 10, 8, 10, 9, 6, 15, 15, 9, 16, 25, 26, 3, 16, 8, 10, 19, 21, 21, 9, 9, 4, 13, 15, 13, 19, 6, 11, 23, 8, 4, 17, 15, 16, 22, 6, 24, 8, 24, 21, 8, 8, 8, 10, 8, 21, 23, 6, 13, 15, 14, 4, 8, 13, 9, 13, 15, 15, 13, 13, 15, 15, 13, 19, 15, 15, 17, 17, 19, 20, 21, 11, 13, 15, 14, 28, 26, 26, 25, 16, 19, 11, 24, 24, 10, 10, 24, 22, 8, 8, 24, 6, 17, 19, 16, 25, 26, 27, 14, 15, 15, 20, 11, 11, 6, 13, 20, 9, 8, 8, 21, 6, 11, 16, 5, 26, 26, 27, 15, 20, 9, 18, 9, 6, 13, 11, 9, 9, 9, 6, 11, 20, 6, 13, 6, 13, 14, 6, 20, 23, 13, 13, 4, 6, 21, 24, 24, 9, 9, 9, 20, 21, 11, 17, 17, 6, 17, 11, 6, 4, 9, 11, 11, 22, 22, 9, 11, 9, 9, 9, 9, 9, 19, 15, 24, 10, 6, 11, 6, 24, 25, 26, 28, 14, 15, 13, 23, 20, 13, 14, 15, 15, 6, 22, 24, 24, 24, 11, 20, 13, 13, 23, 6, 11, 11, 9, 23, 23, 13, 13, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 6, 17, 15, 6, 20, 20, 19, 6, 9, 8, 16, 13, 13, 20, 19, 20, 11, 24, 24, 9, 10, 20, 9, 6, 15, 13, 16, 27, 26, 13, 8, 10, 9, 20, 9, 19, 6, 11, 11, 14, 14, 19, 20, 6, 23, 18, 19, 6, 17, 15, 8, 10, 10, 10, 8, 8, 13, 8, 10, 8, 8, 8, 24, 20, 11, 13, 15, 23, 20, 13, 11, 13, 15, 14, 15, 17, 17, 11, 17, 19, 14, 15, 6, 13, 14, 13, 18, 15, 11, 6, 18, 16, 7, 26, 26, 27, 14, 14, 13, 4, 8, 10, 8, 8, 24, 8, 8, 24, 19, 15, 5, 14, 25, 26, 27, 14, 16, 20, 19, 6, 8, 23, 11, 21, 8, 8, 8, 20, 4, 23, 16, 28, 26, 26, 25, 15, 18, 17, 23, 11, 20, 6, 23, 4, 9, 11, 23, 4, 8, 23, 9, 20, 19, 11, 15, 19, 19, 20, 21, 14, 23, 4, 10, 4, 24, 6, 8, 11, 4, 11, 15, 15, 11, 8, 9, 4, 9, 9, 13, 11, 16, 8, 9, 23, 8, 8, 24, 11, 13, 11, 6, 6, 6, 8, 6, 22, 24, 6, 26, 27, 14, 13, 11, 23, 19, 19, 13, 15, 14, 19, 24, 9, 6, 22, 13, 19, 23, 11, 6, 23, 20, 21, 11, 13, 11, 18, 20, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 11, 19, 22, 8, 9, 23, 20, 11, 21, 22, 9, 20, 19, 11, 11, 19, 11, 8, 11, 6, 22, 20, 8, 8, 19, 19, 17, 26, 27, 15, 20, 9, 21, 15, 13, 15, 19, 11, 15, 13, 18, 20, 8, 23, 9, 8, 20, 17, 13, 8, 22, 8, 10, 8, 8, 10, 4, 22, 24, 8, 10, 8, 9, 20, 13, 15, 13, 4, 14, 15, 15, 15, 14, 14, 11, 13, 15, 6, 6, 14, 14, 20, 6, 13, 15, 13, 20, 13, 11, 9, 20, 24, 16, 27, 26, 26, 25, 14, 19, 20, 8, 10, 8, 10, 10, 22, 8, 4, 14, 19, 13, 13, 7, 28, 28, 19, 8, 24, 11, 13, 9, 9, 9, 13, 20, 8, 23, 9, 6, 16, 7, 26, 26, 27, 14, 5, 17, 13, 9, 9, 19, 11, 4, 9, 23, 23, 6, 6, 11, 13, 24, 21, 10, 10, 9, 19, 13, 20, 13, 13, 21, 23, 9, 9, 13, 24, 6, 9, 11, 15, 22, 24, 22, 22, 20, 4, 8, 6, 15, 13, 8, 8, 8, 6, 21, 20, 6, 4, 11, 4, 8, 8, 11, 4, 4, 6, 24, 15, 27, 26, 17, 19, 20, 13, 13, 11, 4, 24, 19, 15, 14, 6, 11, 11, 21, 23, 20, 20, 20, 13, 20, 20, 20, 13, 21, 11, 16, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 23, 24, 24, 8, 8, 9, 9, 9, 6, 8, 22, 19, 17, 9, 9, 13, 19, 20, 20, 11, 9, 8, 8, 24, 23, 15, 25, 26, 28, 15, 15, 19, 15, 11, 9, 13, 15, 18, 6, 11, 9, 8, 8, 8, 23, 23, 21, 19, 17, 10, 8, 16, 24, 10, 10, 10, 8, 20, 21, 8, 10, 8, 22, 21, 17, 19, 20, 15, 15, 14, 15, 15, 14, 11, 19, 14, 11, 6, 13, 15, 11, 8, 23, 20, 23, 15, 13, 21, 23, 22, 6, 11, 22, 4, 26, 26, 26, 11, 21, 22, 22, 22, 10, 10, 10, 8, 24, 9, 15, 11, 11, 17, 16, 14, 13, 11, 8, 8, 4, 13, 19, 9, 9, 4, 21, 18, 23, 6, 14, 14, 27, 26, 26, 25, 16, 17, 17, 17, 9, 23, 20, 23, 9, 6, 20, 13, 20, 23, 6, 11, 22, 8, 8, 9, 4, 11, 14, 11, 9, 4, 23, 20, 24, 8, 19, 6, 23, 14, 14, 21, 24, 10, 8, 9, 13, 6, 10, 15, 17, 13, 8, 8, 13, 20, 6, 9, 4, 6, 9, 10, 4, 24, 8, 22, 9, 22, 9, 22, 28, 26, 25, 15, 13, 21, 6, 9, 24, 24, 8, 22, 14, 14, 17, 19, 20, 11, 13, 20, 20, 20, 20, 23, 21, 15, 20, 6, 13, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 24, 9, 24, 9, 8, 24, 24, 8, 9, 4, 9, 21, 21, 20, 21, 11, 9, 21, 13, 23, 9, 24, 22, 24, 24, 14, 28, 26, 7, 13, 9, 11, 15, 8, 8, 20, 9, 19, 20, 11, 8, 9, 8, 8, 9, 23, 13, 9, 19, 11, 8, 9, 19, 8, 8, 8, 8, 24, 16, 8, 8, 9, 11, 19, 15, 6, 17, 15, 14, 14, 15, 14, 19, 18, 15, 9, 9, 20, 13, 9, 21, 23, 23, 6, 11, 13, 15, 13, 20, 20, 23, 13, 20, 15, 28, 26, 26, 27, 15, 16, 8, 4, 24, 8, 10, 8, 9, 14, 13, 20, 16, 17, 22, 14, 18, 11, 8, 9, 23, 9, 20, 13, 8, 8, 21, 19, 19, 17, 14, 28, 26, 26, 27, 15, 20, 13, 11, 18, 19, 23, 11, 9, 13, 15, 13, 9, 8, 10, 10, 22, 13, 23, 20, 4, 6, 6, 17, 6, 4, 9, 23, 23, 16, 4, 9, 9, 13, 14, 8, 10, 8, 22, 8, 24, 13, 18, 13, 11, 6, 21, 20, 19, 23, 11, 9, 9, 23, 23, 8, 8, 6, 13, 9, 6, 23, 20, 6, 11, 7, 26, 27, 15, 9, 6, 9, 8, 8, 8, 8, 11, 15, 14, 17, 14, 19, 19, 20, 9, 9, 23, 23, 20, 19, 19, 15, 19, 13, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 8, 9, 8, 24, 8, 9, 8, 8, 24, 8, 20, 8, 23, 19, 18, 20, 20, 23, 14, 15, 18, 19, 22, 8, 5, 16, 26, 27, 15, 22, 8, 11, 19, 11, 4, 11, 6, 6, 11, 23, 6, 6, 13, 11, 9, 20, 11, 20, 13, 23, 13, 9, 6, 18, 8, 10, 10, 24, 22, 6, 6, 13, 13, 14, 17, 17, 15, 15, 15, 14, 17, 11, 13, 11, 9, 9, 19, 23, 13, 9, 23, 20, 9, 9, 20, 23, 19, 19, 23, 6, 20, 20, 19, 21, 16, 27, 26, 26, 28, 16, 8, 8, 4, 9, 22, 23, 6, 15, 6, 20, 22, 6, 6, 25, 3, 15, 24, 13, 9, 9, 9, 11, 21, 11, 21, 15, 18, 16, 25, 26, 26, 26, 4, 22, 15, 9, 4, 11, 14, 15, 21, 13, 13, 23, 23, 6, 5, 8, 8, 18, 21, 20, 8, 19, 21, 8, 9, 13, 15, 23, 6, 8, 9, 19, 6, 19, 14, 9, 10, 10, 8, 10, 10, 4, 8, 21, 15, 21, 21, 14, 21, 23, 6, 23, 6, 23, 20, 8, 8, 9, 6, 20, 8, 4, 8, 15, 19, 17, 14, 27, 26, 5, 22, 4, 8, 4, 8, 8, 24, 6, 13, 14, 15, 11, 13, 17, 13, 23, 20, 6, 20, 13, 11, 14, 13, 15, 22, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 4, 9, 10, 8, 21, 8, 8, 10, 8, 8, 23, 11, 6, 11, 18, 20, 13, 18, 14, 15, 18, 11, 9, 4, 9, 16, 28, 26, 25, 16, 4, 19, 13, 6, 9, 20, 23, 20, 4, 4, 21, 9, 23, 13, 23, 9, 20, 6, 23, 20, 9, 6, 20, 4, 24, 22, 8, 8, 11, 9, 15, 19, 15, 14, 15, 15, 15, 15, 13, 19, 14, 13, 9, 9, 20, 19, 20, 23, 15, 13, 4, 4, 14, 4, 19, 13, 9, 18, 19, 19, 23, 11, 23, 21, 24, 5, 7, 26, 26, 26, 28, 15, 23, 24, 24, 8, 8, 19, 15, 13, 9, 8, 22, 25, 26, 27, 14, 16, 9, 20, 9, 9, 4, 23, 14, 15, 18, 16, 25, 26, 26, 26, 25, 5, 22, 13, 6, 13, 11, 15, 14, 19, 20, 4, 9, 23, 23, 4, 6, 11, 11, 9, 10, 19, 16, 9, 8, 8, 24, 11, 21, 9, 6, 23, 20, 15, 15, 17, 8, 8, 8, 10, 10, 10, 10, 6, 18, 13, 20, 20, 21, 18, 20, 11, 23, 13, 15, 20, 23, 11, 23, 8, 9, 9, 8, 9, 15, 14, 11, 16, 25, 26, 28, 15, 8, 23, 20, 8, 9, 9, 13, 4, 15, 14, 11, 13, 13, 13, 23, 6, 13, 17, 13, 15, 15, 13, 11, 19, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 13, 9, 24, 9, 10, 9, 8, 9, 21, 15, 13, 13, 19, 20, 9, 6, 6, 19, 13, 20, 19, 11, 6, 22, 5, 26, 26, 8, 16, 4, 20, 20, 8, 9, 20, 14, 9, 10, 4, 19, 11, 8, 4, 13, 23, 6, 9, 23, 9, 8, 9, 8, 20, 4, 9, 19, 16, 13, 17, 14, 15, 14, 15, 19, 13, 11, 13, 15, 15, 11, 13, 23, 21, 20, 15, 20, 11, 11, 6, 6, 23, 19, 20, 19, 23, 11, 13, 9, 20, 19, 9, 9, 23, 22, 4, 16, 29, 26, 26, 26, 28, 14, 16, 8, 8, 8, 14, 13, 20, 20, 8, 16, 25, 26, 27, 14, 16, 13, 23, 8, 4, 6, 19, 15, 21, 16, 25, 26, 26, 26, 28, 16, 24, 17, 23, 18, 23, 8, 11, 14, 13, 23, 20, 11, 9, 6, 11, 11, 11, 6, 9, 21, 11, 6, 8, 8, 10, 9, 4, 13, 20, 9, 11, 13, 15, 13, 19, 9, 8, 8, 10, 10, 8, 22, 13, 23, 11, 9, 23, 20, 14, 9, 4, 4, 23, 11, 17, 13, 11, 6, 11, 11, 15, 11, 23, 19, 15, 14, 24, 16, 26, 26, 18, 23, 11, 20, 10, 10, 24, 9, 9, 21, 19, 15, 19, 11, 23, 20, 14, 17, 13, 15, 15, 15, 15, 13, 11, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 4, 15, 9, 23, 20, 23, 23, 23, 21, 15, 22, 8, 24, 24, 9, 9, 8, 23, 22, 8, 8, 9, 15, 7, 16, 12, 26, 28, 16, 13, 6, 9, 9, 21, 9, 23, 19, 23, 4, 6, 23, 9, 8, 6, 13, 11, 9, 8, 22, 9, 8, 9, 9, 20, 18, 17, 15, 15, 15, 21, 6, 15, 14, 13, 13, 11, 21, 19, 21, 20, 4, 17, 13, 15, 13, 11, 11, 13, 9, 8, 9, 22, 9, 15, 13, 4, 6, 11, 6, 9, 21, 23, 8, 6, 13, 6, 13, 14, 29, 26, 26, 26, 27, 17, 16, 24, 17, 15, 8, 8, 24, 19, 14, 25, 26, 27, 15, 24, 18, 8, 9, 6, 15, 21, 16, 13, 28, 26, 26, 26, 28, 14, 15, 14, 23, 23, 23, 23, 4, 21, 21, 20, 9, 19, 19, 20, 9, 20, 18, 9, 6, 15, 19, 8, 8, 10, 10, 8, 22, 6, 20, 18, 11, 6, 18, 8, 8, 14, 6, 4, 8, 9, 9, 16, 9, 4, 9, 11, 11, 8, 8, 22, 16, 9, 23, 20, 8, 4, 20, 9, 9, 24, 13, 17, 13, 14, 17, 11, 14, 9, 16, 28, 26, 25, 15, 6, 8, 4, 9, 4, 4, 21, 11, 20, 15, 15, 20, 20, 19, 20, 19, 14, 19, 11, 21, 14, 19, 13, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 4, 14, 18, 19, 13, 21, 20, 6, 13, 20, 8, 9, 21, 9, 6, 9, 23, 9, 24, 8, 10, 9, 9, 18, 15, 26, 26, 19, 24, 9, 13, 11, 20, 6, 18, 6, 6, 19, 13, 23, 9, 9, 15, 21, 9, 11, 11, 4, 22, 16, 17, 17, 15, 17, 19, 14, 11, 15, 15, 24, 6, 14, 14, 17, 14, 15, 18, 20, 23, 13, 11, 20, 14, 20, 11, 20, 21, 6, 9, 4, 9, 9, 9, 14, 11, 10, 11, 16, 9, 8, 9, 23, 9, 23, 11, 15, 18, 18, 15, 25, 26, 26, 26, 26, 25, 14, 14, 22, 6, 6, 8, 6, 14, 7, 28, 25, 18, 23, 5, 17, 13, 16, 15, 16, 3, 27, 26, 26, 26, 25, 18, 15, 14, 11, 20, 9, 4, 23, 20, 21, 8, 19, 18, 11, 6, 9, 13, 19, 23, 19, 18, 17, 8, 9, 8, 8, 10, 8, 22, 21, 20, 6, 13, 15, 9, 10, 8, 13, 6, 23, 9, 6, 22, 9, 9, 20, 6, 4, 20, 8, 24, 9, 21, 15, 20, 23, 8, 4, 9, 19, 24, 24, 6, 17, 19, 17, 4, 11, 17, 19, 16, 17, 26, 26, 16, 24, 8, 11, 8, 10, 11, 13, 11, 19, 21, 15, 18, 18, 11, 6, 20, 21, 19, 21, 21, 15, 15, 15, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 4, 14, 15, 14, 14, 15, 13, 19, 15, 6, 4, 20, 23, 9, 9, 20, 9, 9, 24, 10, 24, 9, 10, 16, 28, 26, 25, 15, 22, 11, 18, 6, 15, 9, 23, 20, 15, 9, 6, 19, 21, 8, 13, 21, 8, 20, 14, 15, 15, 13, 17, 17, 17, 17, 21, 23, 15, 15, 20, 20, 17, 17, 14, 15, 17, 15, 13, 6, 21, 15, 9, 22, 16, 8, 8, 20, 21, 8, 4, 22, 11, 8, 9, 13, 13, 11, 13, 4, 9, 8, 8, 9, 20, 6, 18, 15, 15, 13, 9, 5, 4, 27, 26, 26, 26, 27, 29, 19, 18, 16, 24, 23, 14, 16, 16, 16, 21, 6, 6, 18, 14, 15, 3, 27, 26, 26, 26, 26, 29, 15, 8, 19, 18, 6, 23, 11, 9, 9, 15, 21, 20, 21, 13, 23, 4, 4, 15, 15, 19, 13, 19, 9, 23, 9, 8, 8, 9, 24, 21, 13, 23, 23, 13, 17, 6, 10, 24, 11, 13, 20, 23, 24, 24, 8, 8, 9, 8, 6, 20, 21, 20, 23, 11, 19, 18, 20, 23, 24, 9, 9, 4, 8, 16, 17, 17, 23, 20, 23, 13, 17, 13, 5, 28, 26, 28, 14, 21, 13, 9, 9, 19, 20, 20, 15, 20, 13, 18, 19, 9, 11, 23, 6, 11, 21, 21, 21, 18, 15, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 15, 13, 11, 17, 15, 20, 18, 15, 15, 19, 17, 6, 11, 20, 20, 9, 11, 9, 22, 22, 8, 5, 10, 26, 27, 16, 8, 13, 17, 13, 9, 18, 11, 4, 8, 13, 4, 8, 17, 15, 20, 20, 20, 21, 23, 13, 17, 17, 6, 9, 23, 23, 9, 8, 23, 21, 13, 9, 20, 15, 14, 11, 15, 13, 11, 23, 20, 15, 6, 24, 22, 8, 8, 10, 23, 8, 8, 8, 24, 9, 6, 9, 20, 19, 19, 16, 9, 8, 8, 9, 9, 23, 21, 23, 11, 14, 11, 23, 9, 16, 15, 28, 26, 26, 26, 26, 26, 28, 25, 8, 15, 14, 14, 24, 15, 14, 16, 24, 29, 28, 27, 26, 26, 26, 26, 27, 6, 14, 13, 11, 13, 15, 23, 9, 4, 17, 14, 14, 15, 11, 9, 20, 23, 9, 19, 18, 20, 13, 18, 11, 11, 23, 8, 8, 24, 9, 9, 21, 19, 9, 16, 6, 6, 16, 9, 21, 6, 6, 4, 15, 24, 4, 4, 4, 9, 9, 20, 19, 15, 6, 6, 6, 6, 23, 23, 20, 6, 4, 4, 13, 22, 6, 11, 17, 23, 21, 23, 24, 17, 11, 24, 16, 27, 26, 4, 16, 4, 9, 22, 20, 13, 20, 18, 19, 21, 21, 20, 15, 6, 9, 20, 23, 23, 11, 19, 21, 22, 4, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 22, 18, 9, 4, 17, 19, 11, 11, 19, 14, 17, 6, 6, 8, 8, 8, 23, 16, 23, 5, 13, 15, 27, 26, 29, 16, 22, 11, 15, 17, 17, 17, 19, 9, 8, 13, 14, 13, 13, 13, 15, 9, 6, 19, 11, 9, 13, 19, 9, 24, 24, 9, 10, 9, 13, 6, 4, 13, 14, 14, 11, 13, 15, 13, 13, 13, 20, 13, 9, 22, 10, 10, 24, 22, 8, 24, 8, 16, 20, 8, 9, 18, 19, 13, 13, 23, 23, 9, 8, 24, 24, 22, 22, 11, 23, 14, 11, 19, 19, 20, 22, 16, 29, 27, 26, 26, 26, 26, 26, 26, 27, 27, 27, 28, 28, 27, 27, 26, 26, 26, 26, 26, 26, 27, 25, 16, 23, 9, 15, 19, 9, 21, 20, 23, 13, 19, 14, 14, 17, 6, 8, 23, 17, 14, 15, 20, 23, 13, 13, 11, 11, 11, 23, 20, 6, 9, 24, 9, 11, 11, 4, 9, 21, 18, 21, 20, 4, 20, 13, 9, 6, 23, 9, 23, 11, 21, 11, 11, 19, 13, 11, 4, 11, 20, 13, 9, 8, 24, 24, 9, 15, 15, 11, 17, 19, 20, 24, 24, 17, 13, 8, 16, 29, 26, 27, 16, 8, 6, 24, 24, 24, 24, 13, 19, 11, 21, 18, 15, 15, 11, 13, 21, 23, 23, 11, 19, 15, 4, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 4, 8, 23, 11, 11, 13, 11, 14, 15, 19, 23, 21, 19, 20, 8, 10, 8, 13, 8, 8, 5, 16, 28, 26, 28, 5, 10, 6, 9, 13, 5, 17, 15, 18, 15, 9, 23, 13, 17, 15, 17, 17, 14, 19, 23, 21, 11, 11, 14, 11, 24, 8, 8, 24, 20, 4, 13, 20, 17, 19, 13, 13, 15, 13, 19, 11, 11, 9, 13, 11, 9, 10, 10, 24, 24, 10, 22, 24, 21, 20, 21, 13, 18, 19, 23, 19, 23, 8, 20, 9, 8, 22, 13, 24, 13, 15, 15, 6, 11, 15, 22, 10, 3, 8, 14, 5, 28, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 27, 29, 5, 5, 23, 9, 23, 20, 13, 20, 6, 18, 21, 19, 20, 11, 19, 13, 15, 20, 20, 15, 14, 9, 8, 20, 19, 6, 11, 18, 15, 19, 9, 9, 8, 4, 4, 19, 11, 20, 21, 20, 9, 11, 18, 6, 21, 13, 6, 11, 21, 18, 13, 23, 9, 9, 9, 6, 21, 11, 19, 23, 6, 6, 21, 24, 24, 9, 9, 17, 17, 13, 17, 19, 8, 8, 8, 13, 19, 4, 20, 15, 28, 26, 28, 16, 24, 8, 8, 8, 22, 19, 17, 23, 6, 15, 23, 13, 15, 23, 13, 18, 20, 23, 11, 18, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 4, 21, 8, 11, 13, 13, 13, 9, 15, 13, 22, 9, 8, 8, 22, 24, 11, 17, 9, 8, 24, 12, 26, 27, 5, 8, 8, 8, 15, 14, 11, 19, 24, 8, 11, 6, 6, 6, 4, 15, 6, 8, 9, 19, 8, 6, 18, 13, 20, 8, 9, 24, 22, 22, 21, 19, 21, 19, 14, 13, 14, 14, 17, 15, 13, 13, 19, 20, 19, 23, 4, 4, 4, 22, 11, 4, 6, 23, 9, 6, 20, 21, 13, 20, 11, 19, 20, 4, 4, 9, 19, 14, 13, 6, 5, 14, 17, 17, 14, 6, 8, 8, 4, 9, 22, 24, 16, 8, 25, 28, 27, 27, 26, 26, 26, 26, 27, 27, 27, 28, 25, 23, 14, 18, 19, 6, 6, 23, 21, 6, 11, 15, 11, 14, 11, 6, 13, 20, 13, 23, 19, 13, 17, 14, 17, 8, 9, 20, 11, 13, 15, 15, 11, 11, 19, 4, 10, 4, 19, 15, 20, 6, 6, 23, 23, 11, 20, 14, 20, 21, 21, 20, 20, 21, 20, 9, 9, 4, 4, 11, 15, 11, 23, 6, 21, 19, 15, 24, 10, 10, 23, 19, 23, 6, 19, 13, 9, 24, 8, 13, 18, 23, 8, 16, 14, 27, 26, 25, 16, 8, 8, 24, 21, 6, 17, 11, 11, 21, 19, 20, 18, 21, 6, 20, 9, 20, 16, 20, 4, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 9, 9, 18, 19, 13, 6, 4, 18, 23, 10, 8, 22, 8, 10, 16, 14, 15, 23, 8, 3, 26, 26, 10, 23, 8, 24, 13, 13, 13, 15, 22, 10, 8, 4, 6, 20, 9, 24, 16, 8, 8, 4, 13, 19, 6, 9, 20, 9, 8, 10, 9, 22, 22, 9, 9, 11, 15, 17, 17, 17, 17, 14, 13, 13, 14, 19, 11, 15, 21, 23, 13, 19, 19, 15, 11, 15, 17, 11, 13, 20, 18, 14, 18, 19, 15, 19, 13, 6, 17, 19, 17, 17, 17, 17, 14, 14, 14, 15, 13, 22, 22, 22, 15, 11, 15, 20, 21, 16, 15, 14, 15, 15, 15, 11, 11, 15, 15, 16, 16, 22, 24, 6, 11, 15, 14, 21, 19, 19, 19, 13, 17, 15, 17, 11, 21, 19, 19, 23, 8, 6, 14, 14, 11, 11, 19, 20, 8, 6, 15, 13, 23, 23, 9, 9, 22, 11, 16, 9, 20, 6, 11, 9, 9, 23, 18, 11, 6, 19, 19, 11, 9, 11, 6, 23, 13, 6, 9, 19, 11, 6, 11, 23, 20, 15, 21, 9, 24, 10, 8, 23, 23, 23, 8, 18, 11, 4, 9, 22, 17, 14, 23, 8, 6, 16, 5, 26, 26, 10, 22, 5, 22, 24, 6, 19, 13, 23, 6, 19, 13, 13, 15, 13, 23, 9, 20, 23, 6, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 10, 22, 16, 15, 17, 11, 16, 8, 10, 24, 4, 4, 11, 17, 23, 23, 11, 14, 11, 26, 26, 29, 16, 8, 9, 13, 15, 11, 20, 14, 15, 4, 9, 6, 9, 19, 24, 24, 24, 9, 22, 21, 23, 23, 21, 11, 19, 19, 8, 11, 18, 18, 13, 9, 17, 14, 15, 15, 17, 6, 6, 6, 15, 17, 14, 19, 9, 21, 8, 9, 20, 21, 23, 20, 19, 14, 21, 11, 6, 15, 19, 14, 17, 14, 15, 11, 15, 15, 15, 11, 6, 4, 18, 14, 15, 6, 15, 13, 8, 8, 8, 17, 20, 23, 18, 6, 9, 9, 11, 19, 24, 11, 18, 14, 22, 17, 21, 8, 8, 8, 6, 24, 8, 23, 13, 14, 14, 11, 13, 19, 15, 17, 14, 15, 15, 20, 13, 23, 11, 19, 15, 15, 20, 13, 19, 21, 20, 19, 18, 6, 23, 23, 9, 6, 11, 14, 6, 4, 13, 13, 23, 8, 4, 9, 19, 20, 17, 13, 15, 17, 11, 11, 23, 9, 11, 13, 17, 9, 4, 9, 15, 11, 22, 9, 9, 8, 9, 20, 20, 9, 9, 8, 20, 23, 18, 20, 23, 8, 6, 21, 19, 11, 24, 8, 16, 29, 26, 26, 4, 16, 9, 6, 11, 18, 21, 6, 6, 11, 13, 23, 11, 15, 21, 19, 19, 11, 9, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 18, 22, 4, 11, 15, 15, 11, 10, 10, 10, 9, 11, 13, 24, 21, 18, 15, 7, 26, 26, 25, 16, 8, 4, 21, 13, 17, 21, 22, 11, 15, 6, 8, 9, 4, 9, 13, 10, 8, 10, 9, 21, 6, 8, 8, 13, 23, 9, 21, 18, 9, 9, 6, 11, 14, 15, 15, 15, 8, 10, 8, 10, 13, 14, 10, 17, 18, 9, 8, 8, 20, 23, 8, 4, 15, 20, 20, 9, 11, 21, 23, 17, 6, 11, 13, 8, 13, 14, 23, 9, 6, 9, 6, 15, 14, 13, 22, 15, 9, 9, 11, 15, 11, 19, 14, 14, 21, 20, 20, 19, 22, 13, 4, 25, 25, 22, 8, 23, 4, 4, 4, 4, 8, 8, 11, 19, 20, 13, 11, 13, 13, 17, 13, 14, 18, 9, 19, 15, 15, 11, 21, 21, 11, 18, 15, 19, 11, 20, 13, 6, 20, 15, 18, 13, 18, 11, 19, 18, 11, 13, 23, 9, 20, 18, 15, 19, 11, 13, 17, 14, 17, 17, 23, 18, 13, 13, 15, 6, 9, 11, 19, 11, 8, 4, 9, 11, 6, 21, 20, 6, 6, 23, 20, 19, 21, 13, 6, 4, 23, 9, 21, 9, 8, 24, 19, 14, 25, 26, 26, 10, 16, 23, 13, 11, 19, 23, 6, 9, 23, 21, 13, 18, 14, 15, 21, 11, 6, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 22, 8, 24, 19, 17, 14, 15, 4, 10, 10, 24, 15, 6, 8, 8, 16, 5, 26, 26, 12, 16, 23, 11, 18, 21, 13, 22, 22, 8, 23, 23, 8, 24, 9, 8, 11, 6, 22, 8, 3, 8, 8, 6, 21, 9, 4, 19, 19, 15, 11, 4, 6, 11, 14, 14, 14, 15, 24, 8, 8, 8, 22, 13, 24, 22, 11, 15, 9, 8, 9, 20, 9, 11, 18, 14, 23, 19, 8, 9, 8, 9, 22, 9, 11, 13, 15, 18, 19, 6, 20, 23, 9, 23, 15, 17, 19, 24, 11, 23, 8, 21, 11, 23, 14, 14, 15, 20, 13, 13, 15, 22, 16, 12, 26, 27, 14, 16, 20, 4, 10, 24, 9, 9, 20, 19, 11, 4, 9, 14, 14, 6, 13, 6, 14, 19, 21, 14, 18, 23, 18, 11, 23, 14, 20, 6, 20, 11, 21, 20, 20, 21, 6, 9, 21, 24, 10, 10, 22, 21, 18, 13, 20, 13, 9, 6, 23, 24, 9, 9, 15, 17, 11, 21, 23, 13, 20, 9, 20, 23, 9, 8, 13, 24, 22, 24, 11, 13, 13, 14, 15, 21, 15, 18, 18, 13, 19, 20, 6, 13, 11, 18, 11, 8, 22, 13, 6, 14, 25, 26, 26, 4, 16, 24, 11, 21, 6, 23, 11, 11, 15, 21, 11, 21, 15, 21, 23, 6, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 8, 9, 22, 9, 17, 15, 14, 15, 15, 19, 13, 4, 23, 8, 5, 29, 26, 26, 25, 14, 6, 17, 18, 20, 4, 21, 21, 8, 10, 23, 9, 10, 24, 24, 13, 24, 4, 22, 8, 10, 8, 10, 10, 13, 15, 13, 18, 18, 6, 23, 21, 23, 13, 15, 14, 14, 6, 5, 5, 8, 24, 22, 24, 10, 22, 15, 19, 22, 9, 19, 11, 13, 15, 14, 13, 13, 6, 24, 22, 10, 8, 8, 8, 22, 22, 22, 13, 15, 20, 11, 23, 23, 13, 15, 13, 6, 22, 19, 13, 9, 13, 6, 15, 15, 23, 11, 23, 23, 19, 11, 8, 5, 25, 26, 27, 16, 5, 13, 16, 9, 9, 23, 23, 18, 11, 11, 18, 19, 13, 19, 15, 13, 15, 13, 19, 14, 19, 9, 18, 23, 13, 15, 15, 20, 8, 19, 14, 15, 4, 4, 4, 9, 11, 23, 8, 24, 24, 8, 19, 15, 15, 13, 6, 23, 6, 8, 8, 10, 8, 19, 15, 13, 23, 23, 20, 9, 8, 8, 8, 10, 10, 20, 9, 4, 4, 6, 17, 11, 15, 15, 21, 23, 23, 11, 23, 13, 11, 21, 15, 9, 18, 16, 8, 22, 8, 6, 17, 14, 25, 26, 26, 29, 16, 20, 13, 19, 19, 19, 21, 21, 15, 21, 20, 15, 13, 19, 15, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 22, 15, 19, 11, 6, 13, 15, 6, 20, 16, 8, 8, 9, 16, 25, 26, 26, 25, 15, 6, 15, 14, 8, 8, 6, 16, 8, 8, 8, 6, 20, 9, 4, 11, 5, 9, 8, 6, 11, 9, 10, 10, 8, 22, 22, 23, 13, 6, 13, 19, 21, 13, 19, 14, 15, 13, 13, 13, 6, 19, 19, 6, 9, 9, 23, 17, 14, 17, 19, 19, 18, 21, 19, 21, 9, 21, 4, 24, 8, 8, 8, 4, 4, 24, 9, 17, 13, 15, 17, 23, 9, 11, 13, 19, 13, 9, 23, 13, 15, 14, 13, 13, 19, 20, 9, 11, 17, 15, 22, 5, 4, 5, 25, 26, 26, 16, 8, 10, 16, 21, 4, 4, 21, 21, 11, 11, 18, 13, 8, 9, 13, 11, 18, 15, 21, 15, 21, 21, 13, 11, 15, 15, 13, 14, 17, 15, 19, 13, 8, 9, 9, 20, 19, 20, 24, 9, 24, 9, 6, 18, 19, 23, 8, 23, 5, 5, 13, 6, 13, 13, 21, 11, 20, 23, 11, 20, 8, 10, 8, 24, 8, 8, 6, 9, 9, 13, 13, 13, 21, 21, 15, 9, 11, 6, 9, 11, 9, 15, 19, 11, 9, 20, 9, 8, 21, 8, 6, 21, 15, 25, 26, 26, 25, 14, 14, 15, 11, 20, 20, 20, 15, 11, 13, 6, 15, 14, 19, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 22, 20, 9, 20, 6, 16, 15, 13, 11, 4, 22, 16, 5, 27, 26, 26, 4, 15, 21, 21, 6, 4, 23, 9, 11, 22, 8, 8, 9, 16, 15, 13, 9, 4, 9, 24, 8, 11, 4, 22, 8, 24, 9, 8, 4, 19, 13, 10, 9, 13, 11, 14, 14, 15, 6, 13, 23, 11, 18, 18, 11, 20, 9, 20, 21, 11, 14, 14, 14, 19, 18, 19, 19, 23, 23, 8, 6, 24, 8, 8, 8, 10, 9, 6, 9, 11, 11, 11, 17, 21, 9, 6, 17, 15, 9, 9, 11, 11, 11, 14, 14, 13, 21, 13, 23, 17, 15, 15, 9, 10, 9, 24, 4, 28, 12, 22, 8, 8, 10, 22, 17, 11, 19, 9, 9, 21, 9, 6, 21, 23, 4, 19, 19, 15, 21, 15, 19, 15, 20, 13, 20, 9, 13, 19, 17, 19, 19, 20, 19, 13, 20, 20, 9, 6, 24, 6, 4, 4, 20, 13, 13, 9, 4, 9, 8, 13, 18, 20, 20, 11, 20, 4, 21, 13, 9, 23, 8, 9, 9, 9, 9, 9, 6, 9, 13, 9, 20, 21, 20, 19, 18, 13, 19, 20, 23, 20, 20, 21, 21, 13, 4, 13, 11, 23, 20, 8, 9, 11, 13, 18, 4, 26, 26, 27, 16, 14, 18, 11, 11, 23, 9, 19, 13, 6, 15, 14, 19, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 9, 8, 23, 8, 23, 4, 15, 19, 20, 16, 16, 29, 26, 26, 27, 16, 16, 9, 24, 9, 9, 9, 9, 11, 18, 23, 9, 9, 19, 23, 4, 15, 11, 9, 8, 6, 6, 9, 6, 16, 22, 10, 10, 24, 24, 9, 24, 4, 10, 4, 14, 14, 14, 24, 24, 9, 8, 20, 21, 11, 13, 23, 9, 20, 9, 13, 15, 15, 14, 19, 18, 21, 11, 23, 23, 9, 15, 13, 24, 9, 8, 4, 11, 9, 4, 4, 13, 13, 6, 20, 23, 11, 13, 19, 9, 6, 20, 13, 15, 14, 19, 15, 18, 23, 20, 15, 17, 11, 22, 10, 9, 8, 24, 16, 16, 24, 10, 10, 10, 24, 19, 14, 8, 4, 6, 9, 9, 8, 9, 11, 19, 15, 19, 15, 19, 15, 15, 19, 20, 20, 19, 21, 22, 4, 15, 11, 11, 6, 23, 20, 15, 13, 23, 20, 11, 9, 4, 9, 15, 6, 11, 11, 6, 13, 21, 23, 9, 23, 23, 21, 20, 19, 21, 11, 6, 20, 20, 20, 13, 22, 13, 16, 19, 20, 20, 9, 11, 19, 13, 21, 13, 18, 15, 21, 11, 21, 14, 18, 15, 13, 21, 15, 15, 13, 21, 20, 13, 14, 19, 15, 15, 15, 27, 26, 26, 25, 15, 16, 14, 19, 21, 18, 15, 13, 17, 19, 11, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 23, 20, 23, 8, 8, 23, 18, 19, 15, 29, 27, 26, 26, 25, 14, 13, 22, 24, 24, 24, 8, 4, 9, 23, 21, 11, 11, 13, 17, 20, 9, 13, 10, 8, 9, 11, 14, 15, 6, 8, 8, 8, 9, 21, 9, 24, 6, 8, 9, 14, 17, 15, 14, 16, 22, 24, 24, 21, 23, 11, 9, 9, 20, 19, 11, 13, 15, 6, 13, 15, 11, 20, 23, 8, 8, 20, 14, 13, 6, 6, 19, 16, 13, 6, 4, 23, 20, 23, 8, 23, 20, 19, 17, 13, 13, 11, 20, 17, 15, 9, 11, 20, 14, 18, 21, 17, 11, 6, 21, 8, 8, 10, 8, 16, 13, 6, 8, 24, 22, 23, 13, 6, 11, 13, 8, 4, 11, 11, 21, 15, 18, 21, 13, 11, 15, 20, 9, 11, 15, 14, 11, 9, 8, 20, 19, 11, 9, 9, 11, 13, 6, 20, 13, 6, 24, 22, 22, 16, 20, 23, 20, 13, 15, 21, 8, 8, 9, 9, 8, 23, 20, 13, 4, 6, 15, 23, 8, 24, 6, 6, 5, 10, 6, 19, 4, 23, 9, 20, 23, 8, 9, 23, 19, 8, 8, 19, 23, 11, 23, 9, 6, 11, 14, 11, 9, 6, 13, 15, 21, 16, 19, 17, 14, 25, 26, 26, 27, 29, 15, 15, 20, 18, 14, 15, 11, 19, 11, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 18, 16, 8, 4, 16, 18, 16, 29, 27, 26, 26, 27, 5, 16, 22, 6, 9, 23, 20, 9, 8, 9, 6, 16, 8, 8, 8, 8, 19, 23, 20, 19, 6, 8, 8, 23, 17, 19, 6, 4, 6, 20, 23, 8, 9, 23, 8, 9, 14, 15, 13, 6, 19, 15, 11, 23, 20, 9, 10, 9, 6, 19, 13, 6, 23, 19, 21, 9, 9, 15, 13, 5, 11, 11, 4, 11, 20, 23, 10, 23, 20, 9, 17, 11, 20, 9, 23, 18, 23, 11, 19, 19, 17, 19, 17, 17, 11, 19, 6, 8, 11, 21, 21, 19, 20, 21, 22, 24, 8, 20, 5, 24, 10, 28, 12, 16, 20, 9, 8, 23, 4, 8, 18, 13, 19, 20, 23, 23, 18, 11, 13, 23, 23, 23, 14, 19, 6, 9, 6, 21, 21, 9, 6, 21, 6, 20, 11, 13, 21, 21, 9, 4, 6, 22, 10, 8, 16, 9, 11, 13, 15, 13, 11, 23, 8, 10, 8, 8, 24, 22, 23, 11, 4, 8, 9, 21, 13, 6, 8, 8, 10, 9, 9, 6, 6, 9, 23, 23, 23, 10, 8, 8, 22, 8, 6, 23, 23, 19, 8, 23, 23, 6, 19, 6, 23, 13, 6, 21, 20, 4, 6, 11, 9, 16, 24, 28, 26, 26, 27, 29, 16, 15, 14, 15, 6, 17, 24, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 22, 23, 16, 14, 5, 12, 27, 26, 26, 27, 3, 16, 20, 22, 8, 10, 22, 6, 4, 13, 9, 9, 13, 16, 4, 8, 24, 8, 9, 23, 9, 23, 13, 22, 22, 9, 17, 13, 21, 13, 9, 11, 19, 23, 23, 20, 8, 14, 14, 13, 15, 4, 23, 17, 19, 4, 8, 9, 11, 9, 4, 11, 9, 23, 8, 18, 20, 9, 4, 13, 11, 11, 13, 13, 8, 23, 9, 21, 20, 18, 8, 6, 6, 9, 8, 8, 23, 19, 9, 11, 15, 14, 19, 14, 14, 19, 15, 14, 23, 8, 9, 19, 6, 13, 21, 23, 19, 11, 4, 13, 4, 24, 12, 26, 27, 15, 9, 9, 19, 11, 11, 13, 20, 9, 10, 6, 13, 9, 9, 23, 8, 9, 23, 13, 15, 11, 19, 20, 8, 4, 9, 20, 9, 23, 9, 6, 21, 20, 6, 9, 20, 8, 9, 23, 18, 16, 9, 6, 17, 6, 9, 11, 17, 23, 21, 10, 8, 9, 9, 23, 9, 13, 11, 23, 24, 9, 11, 9, 24, 24, 9, 22, 8, 9, 11, 9, 23, 20, 8, 4, 10, 24, 8, 21, 20, 4, 18, 13, 9, 13, 6, 6, 11, 14, 21, 21, 9, 13, 11, 4, 4, 20, 19, 13, 13, 14, 4, 27, 26, 26, 27, 25, 17, 14, 15, 15, 16, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 24, 24, 10, 25, 27, 26, 26, 26, 27, 10, 16, 18, 13, 9, 8, 10, 10, 10, 8, 21, 11, 23, 9, 24, 8, 4, 24, 24, 22, 18, 8, 10, 20, 15, 24, 10, 23, 15, 24, 10, 24, 21, 6, 19, 14, 6, 11, 15, 14, 13, 19, 11, 20, 11, 4, 13, 20, 8, 9, 8, 4, 11, 20, 23, 9, 23, 19, 6, 9, 20, 23, 13, 11, 6, 20, 21, 9, 9, 18, 6, 8, 23, 15, 6, 9, 8, 8, 11, 18, 9, 6, 13, 19, 17, 11, 11, 15, 14, 17, 19, 18, 15, 14, 18, 19, 15, 11, 15, 17, 13, 4, 6, 16, 25, 26, 27, 14, 16, 17, 15, 6, 17, 19, 9, 23, 6, 11, 21, 9, 9, 6, 4, 23, 13, 19, 9, 15, 21, 21, 9, 4, 8, 11, 13, 11, 11, 9, 23, 9, 9, 4, 9, 9, 4, 23, 13, 13, 19, 19, 13, 8, 4, 6, 11, 23, 9, 21, 19, 11, 19, 23, 6, 13, 21, 9, 8, 8, 9, 22, 10, 10, 24, 9, 8, 24, 13, 9, 6, 13, 6, 6, 6, 11, 21, 21, 20, 9, 6, 20, 23, 9, 13, 21, 19, 14, 13, 9, 9, 20, 21, 4, 6, 13, 18, 20, 6, 15, 18, 16, 10, 27, 26, 26, 26, 27, 25, 11, 14, 4, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 27, 26, 26, 26, 26, 27, 25, 8, 16, 16, 19, 22, 9, 8, 8, 8, 10, 10, 8, 8, 9, 13, 16, 24, 4, 8, 8, 10, 24, 20, 9, 23, 4, 11, 9, 24, 13, 14, 9, 8, 8, 24, 6, 5, 17, 14, 14, 15, 13, 23, 23, 9, 18, 19, 6, 11, 18, 23, 9, 4, 4, 11, 9, 9, 23, 15, 11, 8, 9, 18, 23, 8, 18, 8, 4, 15, 21, 11, 13, 13, 13, 19, 11, 8, 8, 8, 4, 9, 21, 23, 13, 19, 13, 17, 6, 11, 11, 15, 11, 11, 20, 13, 13, 18, 20, 15, 13, 15, 17, 17, 15, 14, 14, 25, 26, 27, 14, 24, 6, 11, 13, 13, 11, 8, 20, 18, 9, 4, 20, 15, 21, 6, 6, 15, 19, 18, 19, 9, 6, 15, 18, 11, 20, 14, 23, 9, 13, 11, 13, 11, 18, 23, 13, 13, 6, 13, 6, 11, 19, 23, 23, 23, 21, 17, 13, 23, 23, 17, 15, 19, 17, 13, 20, 19, 9, 8, 8, 8, 9, 22, 24, 10, 3, 10, 8, 24, 16, 13, 11, 13, 11, 6, 17, 13, 6, 23, 21, 6, 19, 20, 15, 13, 23, 20, 15, 11, 6, 6, 20, 15, 11, 6, 13, 11, 15, 13, 11, 19, 11, 16, 16, 19, 25, 27, 26, 26, 26, 26, 27, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 2, 26, 27, 27, 12, 8, 24, 16, 8, 23, 17, 21, 8, 9, 8, 21, 8, 10, 10, 10, 10, 10, 9, 16, 21, 9, 4, 8, 8, 21, 20, 8, 10, 10, 24, 24, 10, 13, 15, 13, 15, 23, 9, 24, 23, 4, 15, 15, 15, 13, 18, 23, 13, 18, 6, 18, 8, 6, 15, 21, 23, 18, 16, 4, 9, 19, 15, 13, 9, 21, 9, 8, 8, 24, 16, 6, 19, 14, 19, 6, 15, 14, 8, 24, 8, 10, 10, 4, 8, 23, 19, 20, 20, 6, 15, 11, 23, 18, 13, 13, 15, 6, 17, 13, 9, 20, 11, 13, 14, 15, 17, 24, 16, 14, 7, 25, 25, 15, 19, 11, 15, 13, 11, 23, 13, 6, 9, 11, 11, 9, 20, 20, 6, 13, 15, 15, 20, 11, 4, 9, 23, 15, 21, 20, 4, 23, 19, 9, 8, 19, 13, 13, 6, 18, 19, 6, 9, 8, 9, 9, 19, 9, 4, 13, 17, 13, 11, 13, 15, 17, 11, 17, 6, 17, 15, 19, 19, 13, 20, 9, 20, 18, 4, 8, 8, 24, 22, 15, 21, 19, 18, 19, 6, 15, 11, 6, 13, 19, 14, 15, 20, 11, 23, 13, 11, 20, 13, 9, 21, 13, 20, 13, 6, 9, 20, 20, 15, 21, 15, 13, 11, 9, 15, 18, 14, 11, 29, 28, 27, 26, 2, 1, 1, 1, 1),
		(2, 2, 2, 2, 2, 0, 4, 14, 22, 5, 8, 9, 23, 6, 9, 8, 8, 20, 23, 20, 18, 10, 10, 8, 10, 10, 24, 8, 9, 9, 22, 9, 8, 19, 15, 4, 8, 9, 8, 10, 22, 8, 4, 15, 13, 13, 19, 11, 8, 8, 19, 13, 14, 13, 15, 21, 21, 13, 19, 9, 8, 24, 9, 11, 14, 15, 20, 9, 20, 21, 19, 21, 21, 19, 21, 10, 8, 8, 4, 11, 15, 20, 11, 15, 19, 15, 13, 9, 22, 9, 9, 8, 8, 8, 21, 11, 10, 23, 6, 14, 13, 11, 15, 15, 13, 13, 19, 14, 11, 20, 15, 13, 15, 17, 11, 4, 13, 22, 11, 15, 16, 22, 18, 24, 24, 13, 23, 21, 18, 6, 4, 11, 15, 18, 13, 19, 24, 19, 14, 15, 15, 4, 9, 11, 11, 13, 10, 20, 19, 9, 6, 21, 23, 8, 4, 24, 11, 15, 20, 23, 9, 8, 9, 8, 8, 6, 23, 11, 19, 11, 6, 11, 13, 9, 8, 20, 13, 9, 9, 17, 15, 11, 13, 21, 20, 13, 11, 6, 4, 8, 4, 24, 22, 6, 4, 23, 19, 14, 15, 13, 15, 14, 19, 14, 19, 13, 20, 11, 19, 11, 20, 15, 6, 23, 19, 23, 15, 15, 19, 18, 19, 18, 15, 14, 13, 20, 18, 15, 11, 19, 16, 16, 14, 14, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 18, 14, 20, 6, 13, 19, 23, 8, 23, 6, 23, 21, 19, 11, 6, 8, 10, 10, 9, 10, 8, 8, 10, 8, 16, 18, 8, 6, 9, 22, 24, 8, 9, 16, 24, 6, 17, 9, 23, 13, 9, 9, 13, 17, 17, 17, 19, 19, 23, 4, 11, 15, 20, 10, 10, 23, 6, 13, 14, 21, 18, 20, 13, 21, 19, 6, 19, 23, 11, 23, 22, 10, 8, 19, 20, 9, 11, 15, 15, 11, 22, 9, 24, 9, 8, 22, 20, 20, 10, 8, 20, 13, 11, 6, 15, 14, 14, 15, 15, 15, 15, 13, 20, 19, 9, 13, 4, 21, 8, 8, 22, 6, 15, 15, 15, 13, 8, 10, 6, 13, 11, 9, 6, 13, 18, 23, 19, 18, 19, 18, 19, 11, 14, 17, 23, 13, 11, 6, 23, 6, 23, 9, 14, 20, 8, 13, 8, 4, 8, 20, 11, 23, 13, 20, 10, 8, 24, 8, 21, 6, 21, 15, 20, 9, 11, 23, 8, 8, 9, 21, 11, 4, 9, 21, 13, 23, 8, 20, 11, 8, 21, 21, 6, 4, 9, 9, 11, 13, 11, 20, 15, 15, 14, 14, 19, 13, 11, 17, 9, 9, 11, 8, 6, 9, 11, 9, 10, 6, 11, 11, 23, 11, 6, 9, 9, 20, 14, 21, 11, 15, 19, 19, 13, 6, 6, 11, 14, 8, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 5, 22, 19, 23, 23, 23, 9, 23, 21, 6, 11, 19, 17, 13, 6, 22, 24, 24, 22, 8, 9, 8, 24, 8, 8, 19, 19, 20, 4, 8, 9, 8, 8, 8, 16, 13, 13, 6, 23, 9, 8, 19, 14, 13, 14, 13, 17, 6, 4, 9, 15, 9, 4, 9, 22, 13, 17, 13, 6, 19, 20, 20, 21, 9, 13, 11, 20, 11, 11, 22, 24, 9, 11, 19, 21, 21, 4, 6, 15, 14, 19, 9, 8, 22, 22, 13, 19, 20, 4, 20, 20, 11, 13, 15, 14, 15, 17, 11, 13, 15, 13, 11, 21, 6, 13, 23, 8, 20, 21, 8, 8, 17, 7, 28, 25, 15, 10, 9, 19, 20, 9, 4, 11, 13, 9, 4, 20, 15, 15, 18, 11, 13, 14, 14, 11, 6, 13, 23, 23, 15, 23, 11, 23, 20, 18, 21, 19, 24, 9, 9, 4, 11, 11, 13, 24, 8, 24, 18, 19, 13, 6, 20, 20, 20, 23, 8, 8, 8, 24, 8, 23, 23, 8, 20, 13, 23, 6, 9, 4, 8, 4, 11, 17, 11, 17, 17, 19, 20, 15, 13, 11, 15, 15, 13, 6, 15, 14, 13, 11, 6, 6, 4, 8, 4, 23, 20, 23, 6, 20, 21, 11, 9, 6, 11, 9, 23, 19, 18, 18, 19, 20, 19, 11, 13, 24, 24, 15, 4, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 4, 24, 19, 18, 20, 23, 8, 4, 20, 13, 9, 9, 20, 22, 10, 8, 8, 11, 9, 23, 18, 11, 6, 6, 16, 23, 19, 15, 9, 10, 8, 22, 10, 8, 21, 13, 19, 8, 6, 9, 15, 18, 21, 14, 19, 15, 11, 9, 8, 11, 14, 10, 10, 23, 13, 6, 23, 15, 11, 6, 6, 19, 8, 8, 13, 13, 20, 21, 20, 23, 9, 11, 18, 20, 19, 11, 19, 4, 19, 14, 15, 23, 20, 20, 9, 18, 17, 13, 17, 14, 20, 18, 15, 14, 19, 6, 4, 6, 20, 21, 9, 23, 20, 21, 21, 9, 8, 22, 22, 24, 8, 16, 25, 26, 27, 18, 16, 14, 20, 8, 8, 9, 11, 23, 9, 9, 13, 23, 15, 23, 11, 13, 19, 6, 13, 15, 15, 6, 18, 21, 23, 6, 8, 8, 19, 21, 11, 15, 23, 9, 13, 23, 20, 9, 16, 15, 15, 11, 18, 6, 8, 9, 23, 18, 6, 4, 4, 4, 23, 4, 4, 24, 16, 22, 24, 8, 22, 9, 8, 9, 9, 23, 13, 16, 13, 11, 13, 15, 14, 19, 13, 17, 11, 4, 9, 21, 11, 6, 15, 19, 6, 6, 6, 9, 23, 20, 9, 9, 23, 23, 21, 9, 8, 20, 20, 11, 6, 14, 19, 19, 19, 20, 13, 19, 20, 22, 11, 4, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 11, 22, 11, 19, 15, 21, 9, 9, 20, 19, 4, 6, 13, 24, 9, 10, 24, 6, 11, 18, 20, 9, 9, 22, 4, 10, 23, 8, 23, 22, 24, 8, 9, 19, 15, 15, 15, 11, 11, 18, 15, 20, 18, 11, 19, 13, 14, 19, 18, 17, 6, 6, 16, 19, 6, 10, 13, 21, 15, 13, 21, 23, 6, 23, 14, 19, 20, 9, 23, 9, 11, 21, 11, 8, 23, 21, 19, 17, 11, 13, 14, 15, 20, 9, 19, 15, 19, 15, 15, 19, 11, 19, 19, 13, 9, 20, 6, 20, 6, 11, 4, 6, 13, 19, 15, 20, 8, 9, 24, 24, 13, 16, 25, 26, 27, 14, 22, 17, 18, 11, 9, 23, 4, 9, 9, 20, 6, 20, 15, 20, 6, 6, 15, 20, 23, 23, 13, 11, 11, 11, 13, 13, 22, 13, 6, 23, 20, 6, 18, 4, 8, 6, 6, 13, 19, 20, 21, 19, 15, 6, 6, 11, 19, 6, 9, 23, 9, 8, 6, 4, 4, 9, 8, 9, 16, 9, 9, 23, 23, 9, 23, 23, 6, 13, 15, 13, 19, 19, 4, 8, 18, 15, 6, 9, 11, 20, 11, 11, 9, 15, 18, 21, 13, 6, 8, 20, 8, 23, 21, 9, 19, 21, 8, 9, 21, 20, 9, 15, 23, 18, 13, 19, 13, 13, 13, 22, 6, 4, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 6, 22, 6, 6, 20, 20, 20, 9, 13, 21, 6, 6, 15, 20, 23, 13, 18, 20, 6, 20, 23, 22, 22, 8, 10, 4, 13, 9, 11, 20, 11, 23, 19, 15, 13, 15, 15, 21, 15, 21, 13, 14, 15, 20, 15, 23, 6, 17, 14, 14, 11, 9, 22, 15, 9, 23, 21, 8, 8, 24, 22, 23, 23, 15, 13, 10, 9, 9, 9, 6, 19, 18, 9, 4, 6, 15, 9, 6, 13, 17, 15, 14, 15, 13, 14, 15, 15, 19, 17, 13, 6, 6, 20, 20, 9, 13, 6, 6, 6, 11, 4, 13, 20, 9, 23, 21, 11, 23, 21, 9, 11, 14, 25, 26, 27, 14, 13, 11, 8, 13, 13, 8, 9, 6, 19, 20, 21, 15, 9, 20, 6, 13, 13, 22, 24, 10, 6, 15, 19, 9, 6, 20, 6, 9, 9, 6, 23, 11, 20, 19, 6, 20, 23, 21, 9, 13, 9, 13, 15, 23, 21, 21, 13, 11, 8, 11, 21, 20, 11, 23, 24, 6, 10, 9, 14, 6, 9, 11, 23, 23, 6, 9, 23, 19, 19, 11, 9, 10, 10, 9, 20, 8, 4, 23, 19, 21, 14, 21, 23, 20, 6, 9, 11, 11, 6, 21, 13, 9, 11, 8, 23, 20, 11, 6, 11, 11, 15, 19, 20, 15, 19, 15, 20, 6, 11, 13, 17, 4, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 11, 24, 20, 6, 16, 9, 11, 14, 11, 13, 20, 19, 19, 19, 17, 15, 11, 11, 13, 21, 6, 24, 9, 8, 9, 9, 20, 6, 9, 6, 11, 15, 14, 19, 6, 15, 23, 11, 8, 4, 20, 18, 9, 21, 9, 8, 8, 6, 11, 14, 15, 6, 24, 23, 21, 19, 4, 10, 8, 8, 8, 24, 11, 14, 21, 6, 4, 6, 20, 20, 11, 21, 6, 11, 13, 13, 13, 13, 19, 11, 6, 13, 17, 15, 17, 17, 19, 17, 15, 13, 13, 15, 13, 10, 10, 11, 11, 8, 13, 9, 20, 19, 6, 11, 23, 9, 6, 15, 15, 21, 17, 15, 6, 25, 3, 15, 19, 17, 8, 9, 8, 23, 21, 13, 11, 20, 21, 19, 20, 23, 23, 20, 9, 24, 8, 8, 24, 19, 21, 18, 11, 4, 4, 4, 6, 24, 8, 9, 9, 9, 15, 15, 13, 11, 13, 21, 11, 13, 20, 13, 14, 21, 11, 23, 6, 4, 4, 9, 13, 13, 6, 6, 24, 13, 17, 15, 13, 6, 6, 13, 17, 19, 20, 23, 11, 18, 24, 8, 22, 22, 23, 8, 23, 21, 13, 21, 20, 11, 11, 20, 13, 11, 6, 9, 9, 11, 15, 11, 19, 6, 9, 20, 4, 23, 11, 20, 18, 15, 14, 15, 18, 20, 13, 23, 11, 20, 17, 8, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 6, 8, 9, 6, 11, 19, 23, 11, 19, 22, 8, 24, 24, 16, 19, 11, 11, 9, 13, 4, 6, 24, 10, 10, 10, 9, 15, 20, 6, 6, 19, 19, 20, 11, 23, 15, 20, 8, 10, 24, 22, 23, 20, 20, 8, 9, 20, 23, 9, 20, 19, 13, 18, 18, 18, 6, 4, 8, 22, 24, 24, 13, 11, 13, 8, 18, 20, 21, 21, 6, 13, 13, 15, 21, 9, 9, 18, 9, 10, 22, 8, 14, 13, 15, 14, 20, 6, 13, 15, 13, 19, 14, 22, 8, 23, 13, 13, 9, 17, 9, 20, 20, 6, 13, 13, 13, 11, 11, 15, 15, 15, 11, 15, 16, 24, 17, 15, 19, 18, 8, 8, 21, 18, 19, 13, 13, 17, 19, 21, 9, 8, 20, 20, 23, 8, 6, 21, 15, 8, 23, 19, 11, 8, 20, 23, 8, 8, 4, 9, 11, 20, 13, 19, 11, 13, 6, 21, 9, 20, 13, 15, 19, 13, 19, 20, 20, 9, 9, 19, 21, 9, 8, 11, 9, 9, 19, 9, 9, 23, 11, 11, 20, 11, 23, 20, 23, 21, 13, 11, 18, 15, 19, 18, 9, 19, 14, 23, 6, 23, 13, 20, 13, 21, 23, 20, 23, 18, 23, 11, 20, 13, 19, 9, 6, 13, 17, 13, 14, 14, 11, 17, 17, 9, 17, 13, 19, 17, 4, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 9, 22, 24, 6, 6, 20, 6, 8, 9, 13, 24, 16, 13, 16, 18, 13, 13, 9, 11, 9, 9, 8, 8, 8, 8, 21, 6, 8, 21, 14, 21, 13, 23, 8, 13, 14, 15, 10, 9, 22, 9, 20, 19, 11, 8, 23, 13, 23, 6, 6, 9, 15, 21, 18, 14, 6, 11, 16, 15, 13, 9, 8, 21, 13, 4, 8, 14, 15, 13, 14, 18, 20, 21, 23, 20, 9, 20, 15, 9, 11, 24, 17, 15, 15, 15, 19, 13, 15, 11, 6, 15, 16, 8, 8, 20, 11, 20, 17, 13, 11, 18, 23, 6, 20, 13, 23, 11, 6, 17, 14, 15, 13, 22, 14, 17, 11, 15, 17, 16, 18, 21, 11, 20, 21, 14, 19, 11, 17, 21, 4, 9, 18, 6, 6, 23, 15, 13, 9, 4, 9, 23, 15, 15, 23, 8, 8, 4, 9, 11, 9, 23, 20, 18, 15, 17, 19, 20, 23, 21, 11, 11, 6, 8, 6, 6, 21, 19, 15, 18, 15, 15, 19, 9, 8, 4, 11, 6, 6, 9, 4, 4, 8, 20, 19, 9, 4, 20, 21, 13, 13, 9, 9, 4, 8, 23, 13, 21, 6, 9, 23, 11, 6, 11, 6, 13, 19, 15, 14, 21, 20, 23, 21, 14, 15, 14, 14, 15, 15, 14, 19, 15, 19, 22, 6, 15, 14, 15, 4, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 4, 8, 8, 9, 16, 9, 11, 11, 23, 11, 15, 14, 15, 20, 13, 21, 11, 21, 9, 11, 9, 9, 24, 22, 22, 21, 6, 13, 21, 9, 6, 21, 13, 19, 19, 21, 15, 20, 19, 11, 23, 18, 23, 11, 6, 19, 20, 6, 13, 6, 23, 18, 15, 13, 20, 15, 15, 14, 17, 11, 9, 19, 20, 15, 20, 11, 20, 18, 11, 13, 13, 15, 19, 15, 19, 11, 6, 15, 11, 11, 17, 17, 14, 15, 11, 15, 15, 20, 20, 6, 15, 11, 10, 9, 23, 21, 23, 17, 11, 11, 21, 23, 21, 21, 13, 11, 11, 13, 14, 17, 17, 15, 7, 28, 25, 14, 14, 15, 17, 11, 15, 13, 9, 13, 18, 17, 15, 19, 23, 23, 13, 11, 6, 17, 11, 19, 10, 11, 8, 9, 13, 11, 13, 13, 9, 8, 22, 6, 9, 20, 23, 20, 19, 15, 13, 19, 23, 18, 19, 11, 13, 4, 9, 23, 21, 19, 18, 11, 6, 9, 11, 19, 15, 15, 20, 19, 13, 8, 6, 9, 8, 8, 11, 21, 13, 18, 13, 13, 18, 13, 23, 9, 9, 9, 9, 6, 18, 13, 11, 6, 6, 9, 11, 13, 8, 6, 11, 14, 19, 18, 13, 13, 15, 15, 15, 15, 14, 14, 14, 15, 14, 15, 15, 14, 14, 14, 14, 6, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 4, 8, 8, 24, 11, 9, 6, 18, 19, 11, 13, 14, 15, 11, 6, 21, 20, 15, 13, 9, 9, 23, 20, 13, 6, 19, 13, 11, 4, 8, 6, 6, 15, 19, 19, 20, 15, 17, 19, 11, 17, 13, 6, 21, 21, 11, 11, 11, 19, 11, 13, 6, 13, 21, 9, 19, 14, 15, 15, 17, 15, 13, 20, 6, 11, 21, 9, 20, 15, 13, 18, 14, 18, 13, 20, 6, 8, 19, 17, 11, 5, 15, 14, 14, 13, 9, 20, 14, 8, 6, 14, 9, 8, 6, 4, 9, 9, 19, 17, 13, 20, 8, 6, 11, 23, 20, 16, 14, 15, 17, 17, 16, 25, 26, 27, 14, 14, 15, 19, 13, 17, 19, 21, 20, 11, 11, 17, 19, 20, 20, 17, 11, 13, 17, 11, 20, 8, 23, 9, 6, 11, 6, 6, 13, 15, 20, 9, 9, 24, 6, 9, 6, 8, 17, 15, 4, 9, 15, 15, 15, 19, 20, 11, 23, 18, 20, 9, 9, 11, 11, 11, 20, 13, 21, 23, 8, 21, 23, 13, 21, 21, 18, 15, 13, 21, 20, 11, 11, 9, 15, 13, 20, 13, 11, 13, 21, 23, 21, 19, 21, 11, 9, 4, 23, 11, 9, 9, 19, 13, 9, 11, 19, 14, 14, 14, 14, 14, 14, 14, 14, 15, 19, 11, 13, 14, 14, 14, 6, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 4, 8, 24, 8, 22, 20, 20, 21, 23, 8, 13, 19, 9, 18, 13, 11, 19, 19, 11, 8, 6, 6, 19, 20, 23, 18, 9, 8, 8, 8, 9, 21, 24, 9, 15, 13, 14, 15, 11, 20, 15, 11, 11, 21, 23, 6, 11, 6, 19, 22, 4, 8, 24, 19, 15, 17, 19, 6, 11, 21, 14, 9, 6, 6, 9, 23, 13, 23, 19, 14, 22, 8, 8, 24, 24, 19, 19, 21, 15, 6, 13, 20, 13, 14, 13, 6, 20, 18, 19, 11, 13, 11, 8, 4, 4, 8, 9, 21, 24, 22, 22, 23, 13, 6, 4, 6, 14, 11, 23, 13, 15, 15, 25, 26, 27, 14, 19, 4, 19, 15, 21, 19, 14, 15, 11, 11, 11, 6, 20, 19, 13, 13, 11, 13, 19, 9, 9, 11, 11, 24, 8, 24, 22, 22, 22, 16, 13, 9, 8, 4, 4, 9, 8, 13, 15, 17, 13, 17, 14, 14, 23, 9, 9, 23, 20, 6, 20, 6, 20, 19, 17, 20, 8, 8, 22, 9, 6, 6, 8, 9, 21, 15, 19, 19, 17, 11, 14, 17, 11, 19, 19, 23, 6, 13, 23, 13, 9, 9, 11, 23, 20, 9, 4, 9, 13, 21, 20, 19, 15, 21, 21, 11, 19, 14, 15, 19, 17, 14, 15, 15, 13, 13, 17, 13, 15, 15, 17, 6, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 4, 24, 8, 24, 22, 24, 8, 4, 9, 10, 21, 20, 8, 24, 21, 6, 19, 6, 23, 4, 9, 20, 23, 9, 23, 22, 8, 8, 8, 10, 24, 8, 8, 4, 19, 13, 19, 15, 6, 19, 13, 18, 21, 13, 9, 11, 9, 19, 15, 9, 9, 21, 24, 9, 20, 18, 9, 4, 10, 23, 9, 11, 14, 11, 9, 4, 20, 11, 18, 13, 6, 10, 8, 22, 22, 24, 11, 15, 14, 14, 23, 11, 19, 18, 14, 13, 18, 23, 14, 19, 17, 22, 24, 24, 6, 23, 23, 8, 24, 9, 8, 8, 11, 6, 19, 21, 11, 4, 9, 19, 15, 18, 25, 26, 27, 14, 15, 11, 21, 20, 9, 13, 19, 17, 19, 11, 23, 21, 20, 13, 13, 15, 11, 13, 23, 8, 11, 11, 13, 8, 22, 22, 24, 8, 10, 10, 6, 22, 10, 4, 9, 9, 24, 13, 6, 14, 15, 6, 17, 15, 23, 8, 6, 9, 21, 9, 6, 23, 15, 13, 6, 23, 24, 8, 24, 22, 15, 19, 9, 23, 21, 15, 20, 23, 9, 23, 11, 6, 15, 19, 20, 13, 9, 23, 23, 13, 9, 8, 11, 11, 13, 19, 21, 23, 6, 19, 23, 21, 15, 9, 8, 9, 13, 15, 13, 11, 17, 14, 15, 14, 13, 11, 13, 15, 13, 11, 17, 6, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 9, 8, 24, 24, 9, 8, 8, 10, 24, 23, 19, 23, 9, 8, 8, 22, 15, 23, 9, 6, 21, 20, 8, 6, 18, 24, 9, 9, 8, 21, 9, 10, 8, 9, 19, 9, 19, 13, 20, 21, 20, 18, 19, 13, 11, 13, 13, 15, 13, 24, 24, 9, 10, 10, 8, 15, 24, 10, 9, 23, 9, 21, 15, 13, 4, 10, 9, 15, 19, 10, 8, 19, 6, 8, 9, 24, 13, 13, 20, 13, 15, 18, 23, 4, 14, 19, 11, 9, 18, 19, 19, 9, 10, 4, 9, 11, 21, 8, 9, 24, 24, 8, 6, 20, 13, 19, 20, 21, 15, 14, 19, 19, 17, 25, 4, 15, 15, 14, 21, 18, 21, 15, 17, 13, 13, 13, 18, 13, 6, 11, 13, 15, 13, 15, 20, 6, 6, 6, 13, 9, 8, 10, 10, 8, 8, 4, 6, 13, 22, 9, 4, 9, 13, 23, 20, 20, 14, 11, 11, 13, 23, 21, 21, 11, 11, 6, 8, 19, 15, 4, 6, 21, 22, 22, 22, 8, 6, 17, 23, 23, 11, 20, 9, 8, 8, 24, 4, 8, 6, 13, 9, 11, 19, 13, 13, 15, 20, 11, 6, 19, 20, 11, 13, 9, 4, 11, 20, 8, 14, 20, 8, 24, 15, 19, 8, 23, 15, 19, 13, 19, 11, 11, 19, 19, 9, 24, 15, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 17, 8, 8, 8, 8, 8, 8, 8, 24, 21, 23, 23, 4, 8, 8, 16, 11, 13, 8, 19, 6, 4, 6, 11, 11, 24, 9, 9, 21, 21, 8, 24, 8, 20, 20, 9, 23, 20, 15, 9, 21, 18, 19, 13, 13, 13, 9, 21, 11, 22, 24, 10, 4, 10, 8, 8, 16, 20, 18, 23, 20, 23, 8, 10, 21, 19, 6, 20, 9, 8, 8, 24, 19, 24, 8, 11, 17, 17, 21, 20, 19, 21, 20, 21, 21, 19, 19, 11, 21, 13, 17, 21, 8, 10, 9, 23, 23, 10, 24, 8, 8, 23, 13, 4, 11, 6, 23, 23, 13, 19, 15, 17, 22, 22, 22, 14, 19, 15, 18, 11, 14, 15, 13, 14, 17, 19, 14, 15, 13, 14, 19, 13, 19, 14, 15, 19, 19, 11, 11, 9, 10, 8, 9, 24, 24, 8, 9, 4, 6, 19, 24, 6, 4, 9, 8, 4, 9, 15, 15, 13, 15, 20, 21, 18, 19, 13, 19, 13, 13, 19, 13, 24, 8, 10, 10, 8, 9, 17, 15, 13, 6, 4, 8, 8, 22, 24, 8, 21, 16, 9, 6, 23, 13, 21, 6, 20, 9, 11, 9, 11, 18, 6, 8, 11, 13, 4, 6, 11, 21, 21, 24, 15, 11, 11, 24, 24, 19, 11, 13, 17, 13, 17, 23, 20, 23, 24, 19, 3, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 6, 22, 10, 9, 8, 10, 8, 8, 9, 8, 11, 20, 9, 8, 24, 22, 10, 20, 14, 9, 4, 9, 13, 4, 24, 8, 9, 22, 13, 9, 11, 9, 11, 4, 13, 6, 20, 14, 18, 21, 19, 23, 6, 11, 20, 4, 23, 19, 4, 6, 9, 4, 4, 11, 24, 8, 24, 14, 13, 9, 9, 8, 20, 23, 8, 4, 14, 13, 8, 8, 9, 8, 22, 19, 21, 13, 13, 13, 18, 23, 23, 19, 6, 9, 21, 15, 15, 19, 9, 21, 11, 11, 15, 8, 8, 24, 24, 9, 8, 9, 13, 18, 8, 22, 22, 9, 8, 10, 22, 18, 11, 6, 16, 14, 18, 14, 13, 5, 17, 14, 14, 13, 17, 11, 22, 16, 23, 20, 14, 14, 13, 19, 6, 10, 18, 19, 13, 6, 9, 11, 24, 23, 6, 6, 11, 13, 13, 11, 13, 11, 14, 18, 11, 20, 23, 9, 13, 14, 14, 15, 17, 15, 20, 11, 23, 15, 14, 11, 13, 9, 8, 10, 10, 10, 10, 10, 8, 24, 15, 17, 17, 6, 23, 23, 21, 9, 22, 24, 9, 10, 10, 8, 11, 22, 22, 8, 10, 8, 9, 9, 19, 15, 19, 6, 11, 20, 9, 6, 11, 17, 17, 19, 8, 24, 19, 16, 21, 8, 13, 15, 13, 19, 18, 18, 13, 16, 17, 3, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 4, 8, 8, 24, 9, 8, 10, 24, 8, 8, 19, 19, 9, 9, 22, 8, 8, 23, 21, 23, 9, 24, 4, 4, 24, 4, 11, 9, 9, 9, 8, 11, 6, 23, 19, 23, 14, 20, 21, 11, 23, 8, 21, 11, 4, 23, 15, 6, 9, 11, 24, 24, 6, 22, 8, 4, 6, 15, 11, 15, 8, 23, 23, 4, 8, 11, 15, 19, 20, 9, 24, 8, 10, 20, 14, 17, 17, 19, 13, 11, 13, 15, 9, 8, 4, 21, 18, 14, 13, 21, 13, 9, 13, 14, 9, 9, 8, 24, 6, 21, 15, 22, 9, 8, 10, 10, 10, 8, 21, 8, 5, 13, 29, 27, 28, 14, 17, 13, 19, 14, 15, 19, 11, 11, 22, 22, 23, 6, 15, 11, 9, 14, 20, 21, 21, 6, 13, 8, 10, 10, 3, 10, 6, 11, 20, 19, 20, 23, 11, 23, 13, 21, 15, 20, 9, 8, 9, 14, 14, 15, 17, 15, 21, 15, 18, 14, 13, 21, 19, 9, 9, 22, 21, 24, 9, 24, 22, 15, 14, 23, 18, 19, 8, 23, 9, 20, 24, 8, 8, 10, 8, 10, 4, 6, 21, 22, 8, 8, 9, 11, 20, 13, 23, 6, 6, 20, 16, 11, 17, 14, 15, 4, 9, 24, 15, 23, 20, 23, 13, 15, 19, 11, 19, 18, 15, 23, 11, 10, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 9, 8, 8, 22, 8, 8, 22, 21, 24, 11, 9, 6, 11, 6, 9, 24, 24, 4, 4, 21, 19, 6, 10, 6, 13, 11, 4, 6, 13, 11, 20, 20, 4, 13, 13, 11, 18, 23, 19, 20, 23, 11, 21, 20, 9, 23, 13, 6, 19, 13, 11, 4, 6, 6, 4, 4, 24, 13, 17, 11, 18, 21, 8, 9, 20, 17, 13, 19, 20, 8, 10, 10, 8, 8, 23, 19, 17, 13, 6, 13, 21, 6, 6, 4, 8, 21, 21, 9, 14, 14, 13, 9, 23, 19, 21, 21, 23, 13, 15, 18, 11, 23, 8, 10, 10, 10, 8, 21, 8, 8, 5, 15, 25, 26, 27, 14, 19, 17, 14, 15, 15, 14, 13, 11, 22, 24, 11, 13, 20, 8, 19, 20, 9, 11, 6, 9, 4, 20, 11, 22, 9, 24, 24, 9, 9, 23, 9, 23, 23, 18, 23, 19, 15, 21, 9, 4, 23, 17, 14, 11, 19, 15, 18, 23, 6, 6, 8, 11, 21, 11, 24, 24, 24, 9, 10, 8, 21, 9, 22, 22, 24, 9, 19, 13, 20, 21, 24, 9, 22, 8, 24, 22, 22, 6, 19, 15, 18, 21, 19, 20, 11, 20, 13, 6, 9, 9, 24, 21, 15, 14, 17, 6, 24, 24, 17, 11, 13, 6, 13, 15, 13, 11, 13, 13, 15, 16, 11, 3, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 9, 8, 10, 22, 9, 9, 24, 8, 24, 13, 4, 9, 19, 9, 24, 8, 10, 10, 4, 18, 8, 23, 6, 9, 19, 9, 6, 13, 4, 11, 9, 8, 9, 19, 23, 11, 23, 20, 23, 19, 23, 23, 19, 23, 23, 13, 19, 20, 11, 6, 4, 23, 19, 8, 10, 9, 22, 11, 17, 18, 20, 15, 6, 13, 11, 17, 11, 9, 23, 8, 8, 10, 24, 23, 8, 6, 15, 6, 9, 19, 21, 4, 6, 9, 6, 13, 18, 4, 15, 18, 23, 20, 18, 13, 6, 14, 15, 19, 18, 8, 6, 21, 10, 10, 4, 24, 24, 24, 8, 9, 6, 16, 25, 26, 27, 14, 18, 15, 17, 13, 17, 17, 14, 13, 22, 17, 17, 6, 23, 4, 23, 13, 11, 10, 9, 21, 13, 15, 11, 19, 24, 8, 10, 10, 8, 8, 4, 9, 21, 23, 11, 19, 6, 23, 21, 14, 14, 17, 18, 13, 9, 15, 14, 21, 11, 6, 6, 9, 21, 20, 22, 8, 10, 8, 10, 9, 24, 10, 24, 22, 8, 10, 9, 6, 19, 4, 8, 10, 9, 8, 8, 24, 16, 6, 6, 17, 14, 13, 6, 23, 19, 11, 20, 21, 6, 23, 24, 23, 14, 14, 15, 6, 22, 15, 14, 14, 15, 15, 14, 13, 15, 11, 11, 21, 14, 14, 17, 8, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 4, 8, 8, 6, 24, 21, 10, 10, 8, 22, 9, 11, 13, 19, 9, 10, 10, 8, 22, 8, 22, 4, 18, 15, 4, 10, 22, 10, 8, 8, 4, 22, 24, 6, 6, 8, 20, 4, 4, 17, 11, 13, 16, 9, 24, 9, 11, 24, 24, 9, 6, 21, 9, 8, 8, 21, 21, 21, 13, 11, 13, 18, 19, 11, 6, 6, 8, 8, 9, 4, 23, 13, 23, 23, 4, 9, 22, 20, 13, 20, 23, 8, 9, 21, 17, 21, 21, 13, 13, 15, 23, 18, 23, 17, 17, 14, 15, 13, 9, 6, 19, 9, 9, 9, 6, 23, 9, 20, 9, 23, 6, 16, 25, 26, 27, 17, 16, 17, 13, 17, 6, 13, 14, 14, 17, 15, 19, 11, 23, 20, 9, 9, 9, 13, 11, 23, 24, 24, 6, 9, 9, 9, 8, 10, 8, 8, 8, 21, 13, 6, 6, 6, 6, 13, 15, 14, 15, 19, 18, 18, 21, 6, 15, 19, 9, 6, 6, 9, 6, 4, 8, 24, 24, 10, 9, 9, 10, 8, 8, 22, 10, 8, 8, 20, 6, 23, 23, 6, 13, 8, 8, 8, 24, 24, 13, 6, 6, 19, 23, 8, 23, 6, 11, 11, 11, 8, 8, 20, 18, 23, 14, 11, 13, 22, 6, 18, 20, 15, 14, 21, 18, 15, 15, 15, 6, 18, 13, 8, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 13, 22, 20, 6, 11, 21, 8, 8, 22, 22, 24, 6, 15, 14, 8, 24, 24, 21, 10, 10, 9, 6, 9, 23, 6, 24, 9, 9, 8, 8, 22, 22, 8, 20, 6, 8, 20, 9, 19, 15, 11, 6, 9, 10, 8, 6, 13, 8, 24, 9, 11, 11, 4, 9, 15, 14, 13, 23, 13, 9, 20, 21, 6, 20, 23, 6, 6, 9, 24, 8, 6, 13, 13, 10, 10, 13, 6, 20, 20, 23, 4, 10, 8, 20, 14, 20, 21, 19, 17, 11, 15, 13, 6, 15, 14, 6, 21, 15, 23, 18, 21, 23, 20, 20, 6, 8, 23, 8, 23, 24, 11, 22, 11, 25, 4, 19, 14, 15, 15, 11, 20, 15, 11, 17, 17, 14, 23, 11, 21, 13, 6, 9, 9, 6, 19, 21, 10, 10, 4, 9, 9, 9, 22, 22, 22, 9, 22, 11, 23, 19, 15, 15, 15, 13, 6, 20, 9, 19, 21, 20, 20, 23, 19, 14, 19, 21, 24, 4, 9, 10, 10, 10, 8, 19, 24, 10, 8, 9, 4, 11, 9, 9, 22, 24, 4, 9, 20, 20, 11, 8, 8, 24, 22, 9, 11, 9, 8, 9, 18, 21, 6, 6, 11, 9, 13, 20, 23, 13, 21, 20, 17, 14, 11, 8, 6, 14, 20, 4, 23, 9, 19, 14, 19, 13, 6, 14, 13, 3, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 9, 24, 6, 22, 4, 8, 21, 8, 8, 22, 8, 11, 14, 13, 6, 8, 16, 8, 10, 10, 8, 20, 10, 20, 4, 22, 22, 8, 8, 9, 8, 10, 10, 19, 13, 13, 19, 18, 8, 8, 24, 8, 9, 8, 10, 13, 11, 8, 8, 9, 19, 6, 11, 19, 14, 13, 20, 9, 21, 8, 6, 18, 4, 23, 19, 4, 4, 9, 11, 6, 13, 23, 9, 9, 9, 13, 11, 4, 11, 15, 23, 8, 8, 9, 14, 9, 22, 15, 15, 13, 19, 14, 13, 11, 19, 14, 23, 23, 15, 15, 11, 23, 23, 20, 4, 4, 23, 11, 21, 22, 13, 15, 16, 16, 18, 14, 11, 16, 8, 8, 22, 9, 9, 17, 14, 6, 9, 6, 18, 20, 19, 21, 23, 6, 6, 19, 8, 10, 10, 4, 22, 9, 8, 15, 15, 9, 20, 20, 22, 22, 24, 24, 22, 8, 9, 10, 24, 15, 19, 4, 23, 11, 8, 13, 14, 11, 13, 11, 11, 10, 8, 10, 8, 8, 8, 9, 9, 9, 9, 24, 16, 24, 8, 10, 8, 10, 8, 20, 23, 9, 24, 22, 9, 4, 9, 9, 6, 9, 9, 15, 20, 6, 9, 8, 9, 14, 14, 14, 15, 13, 17, 14, 16, 9, 20, 15, 8, 4, 23, 19, 19, 15, 9, 9, 23, 15, 6, 3, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 10, 10, 9, 6, 9, 9, 24, 8, 8, 24, 24, 6, 6, 9, 6, 22, 10, 10, 8, 24, 8, 4, 11, 19, 8, 23, 16, 22, 8, 8, 8, 8, 22, 14, 11, 20, 13, 10, 3, 10, 22, 9, 9, 8, 9, 19, 4, 8, 10, 20, 6, 6, 15, 14, 20, 20, 9, 9, 11, 20, 20, 20, 6, 9, 8, 11, 6, 6, 11, 21, 9, 4, 8, 6, 19, 15, 10, 8, 6, 23, 13, 21, 9, 16, 15, 21, 24, 13, 14, 17, 11, 14, 21, 11, 15, 8, 9, 23, 18, 15, 11, 11, 21, 11, 20, 15, 15, 17, 13, 22, 6, 11, 20, 22, 14, 11, 13, 24, 8, 24, 8, 9, 16, 24, 11, 19, 9, 14, 11, 4, 23, 4, 6, 13, 13, 20, 22, 24, 8, 9, 22, 9, 4, 6, 13, 14, 14, 21, 10, 10, 24, 22, 10, 8, 24, 10, 8, 16, 20, 9, 19, 21, 10, 8, 20, 11, 9, 8, 24, 8, 24, 21, 21, 9, 9, 8, 24, 8, 10, 4, 19, 8, 10, 10, 8, 8, 10, 11, 21, 16, 8, 9, 9, 23, 6, 9, 8, 9, 9, 9, 13, 13, 6, 9, 13, 13, 14, 17, 15, 17, 13, 17, 13, 22, 15, 6, 6, 11, 15, 21, 9, 21, 20, 11, 19, 11, 6, 3, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 4, 8, 22, 24, 8, 8, 9, 23, 20, 8, 8, 8, 8, 24, 24, 24, 10, 8, 24, 8, 10, 9, 14, 9, 20, 22, 8, 21, 16, 23, 9, 9, 11, 15, 21, 23, 4, 10, 10, 10, 22, 11, 20, 9, 13, 8, 3, 8, 24, 17, 6, 19, 15, 23, 24, 24, 9, 8, 23, 13, 18, 8, 10, 9, 10, 9, 19, 11, 15, 9, 8, 10, 8, 16, 19, 19, 9, 6, 20, 23, 19, 14, 13, 15, 23, 18, 13, 13, 14, 19, 13, 23, 15, 15, 19, 9, 23, 13, 21, 13, 15, 15, 23, 20, 19, 15, 16, 9, 10, 8, 8, 24, 29, 27, 28, 19, 18, 5, 23, 11, 6, 24, 22, 9, 10, 19, 15, 13, 24, 6, 23, 8, 9, 8, 9, 13, 11, 15, 13, 6, 6, 9, 13, 19, 13, 20, 11, 21, 6, 9, 22, 8, 8, 24, 9, 24, 9, 23, 11, 21, 22, 9, 9, 23, 4, 21, 13, 9, 8, 13, 22, 24, 9, 22, 24, 8, 10, 9, 11, 21, 11, 4, 8, 10, 8, 24, 6, 19, 9, 9, 9, 11, 9, 23, 23, 9, 9, 8, 6, 6, 20, 18, 13, 18, 13, 11, 15, 13, 11, 15, 11, 21, 21, 23, 20, 21, 15, 14, 9, 11, 20, 19, 18, 6, 11, 19, 15, 9, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 17, 16, 16, 8, 4, 8, 8, 20, 18, 8, 10, 8, 8, 21, 10, 8, 8, 24, 9, 8, 9, 4, 21, 21, 14, 22, 8, 9, 9, 23, 8, 11, 19, 16, 8, 8, 9, 8, 10, 8, 9, 18, 9, 4, 13, 10, 10, 10, 15, 11, 23, 21, 11, 8, 8, 8, 8, 9, 11, 11, 15, 10, 8, 24, 10, 8, 6, 14, 11, 9, 8, 8, 9, 20, 11, 6, 6, 21, 21, 11, 23, 13, 14, 15, 9, 20, 19, 17, 14, 18, 11, 11, 15, 14, 20, 11, 21, 23, 21, 19, 20, 21, 21, 6, 9, 8, 8, 9, 9, 23, 4, 8, 25, 26, 27, 14, 24, 22, 18, 11, 13, 23, 9, 10, 10, 11, 14, 9, 10, 9, 19, 11, 4, 23, 6, 11, 9, 6, 13, 14, 15, 13, 20, 9, 9, 9, 4, 8, 18, 19, 24, 9, 8, 22, 23, 8, 23, 23, 13, 24, 8, 10, 11, 20, 9, 23, 19, 15, 20, 9, 8, 8, 10, 8, 8, 10, 8, 4, 19, 19, 19, 23, 24, 8, 9, 24, 9, 20, 9, 9, 23, 20, 6, 23, 9, 9, 6, 6, 6, 11, 19, 19, 18, 21, 11, 19, 11, 11, 14, 11, 23, 19, 18, 6, 15, 21, 14, 19, 9, 19, 6, 13, 11, 23, 18, 19, 14, 4, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 6, 24, 18, 20, 20, 6, 8, 23, 21, 9, 24, 24, 9, 9, 8, 10, 22, 8, 10, 10, 9, 20, 15, 14, 11, 22, 8, 8, 10, 4, 13, 15, 15, 24, 8, 8, 8, 8, 8, 24, 6, 19, 10, 8, 9, 10, 4, 13, 13, 11, 21, 21, 10, 10, 8, 8, 8, 23, 6, 9, 6, 10, 24, 3, 24, 20, 13, 11, 11, 11, 9, 6, 21, 9, 20, 23, 20, 19, 15, 23, 6, 11, 14, 15, 21, 23, 14, 15, 14, 23, 23, 13, 21, 15, 18, 15, 13, 20, 14, 23, 8, 9, 20, 13, 23, 8, 8, 8, 24, 20, 8, 16, 25, 26, 27, 15, 13, 15, 20, 20, 9, 8, 10, 8, 24, 21, 15, 6, 9, 4, 13, 21, 8, 6, 11, 13, 11, 23, 8, 11, 18, 11, 23, 20, 13, 4, 4, 23, 23, 13, 13, 8, 19, 15, 23, 9, 23, 9, 17, 10, 8, 24, 15, 20, 9, 9, 6, 15, 19, 8, 8, 8, 9, 8, 8, 8, 10, 9, 13, 4, 4, 15, 13, 24, 24, 6, 20, 13, 23, 23, 11, 6, 9, 20, 9, 4, 4, 23, 13, 19, 19, 11, 14, 13, 18, 15, 13, 15, 14, 6, 6, 9, 21, 15, 14, 11, 6, 15, 19, 21, 9, 9, 21, 15, 15, 24, 6, 4, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 10, 23, 23, 13, 11, 13, 13, 15, 11, 13, 4, 22, 19, 8, 4, 8, 24, 10, 8, 8, 24, 22, 23, 19, 13, 9, 8, 24, 8, 9, 23, 19, 13, 17, 8, 8, 10, 8, 24, 22, 9, 8, 6, 9, 11, 20, 24, 19, 19, 6, 22, 22, 8, 10, 10, 8, 9, 24, 6, 23, 4, 13, 9, 9, 4, 24, 15, 6, 9, 23, 11, 6, 19, 17, 13, 15, 11, 13, 20, 23, 13, 21, 17, 14, 20, 20, 19, 6, 17, 17, 11, 15, 19, 14, 14, 14, 18, 9, 11, 15, 23, 20, 23, 9, 6, 13, 23, 8, 9, 9, 8, 8, 14, 25, 26, 27, 15, 11, 11, 11, 20, 4, 4, 8, 24, 22, 19, 13, 11, 22, 16, 20, 9, 18, 13, 6, 23, 9, 4, 8, 4, 9, 19, 9, 6, 9, 13, 19, 20, 9, 4, 6, 15, 17, 6, 6, 13, 19, 15, 11, 10, 10, 8, 9, 11, 8, 4, 20, 15, 20, 18, 8, 8, 10, 8, 8, 10, 4, 19, 8, 4, 8, 16, 11, 6, 6, 6, 11, 13, 11, 21, 13, 6, 4, 9, 11, 13, 21, 19, 13, 13, 21, 14, 13, 13, 19, 13, 14, 15, 9, 17, 9, 9, 13, 19, 9, 18, 19, 15, 23, 19, 9, 11, 15, 20, 9, 18, 17, 4, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 24, 9, 8, 4, 9, 16, 6, 11, 17, 19, 18, 20, 20, 13, 19, 9, 4, 22, 22, 8, 10, 22, 9, 8, 16, 23, 21, 20, 6, 15, 16, 4, 13, 8, 8, 10, 6, 9, 24, 22, 8, 11, 11, 11, 17, 11, 21, 19, 11, 9, 20, 9, 6, 9, 4, 4, 4, 23, 8, 23, 6, 9, 4, 6, 24, 6, 23, 11, 21, 15, 14, 13, 23, 13, 17, 6, 22, 18, 11, 9, 17, 15, 17, 11, 17, 19, 13, 15, 17, 15, 16, 19, 15, 21, 18, 19, 15, 15, 20, 23, 4, 4, 9, 19, 4, 9, 9, 23, 23, 4, 16, 23, 17, 7, 13, 20, 10, 6, 13, 9, 4, 10, 9, 8, 11, 17, 6, 13, 15, 14, 15, 20, 11, 13, 22, 9, 4, 10, 8, 8, 8, 11, 15, 20, 4, 6, 9, 8, 11, 11, 17, 14, 17, 11, 11, 9, 15, 19, 11, 10, 8, 8, 10, 10, 13, 13, 9, 11, 20, 6, 16, 8, 10, 8, 8, 8, 17, 6, 8, 22, 8, 8, 9, 6, 20, 9, 23, 6, 9, 6, 13, 15, 15, 14, 18, 19, 20, 9, 8, 11, 15, 11, 8, 13, 15, 13, 19, 13, 13, 15, 18, 6, 11, 19, 10, 9, 15, 19, 6, 6, 15, 13, 21, 9, 10, 8, 17, 8, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 7, 24, 6, 4, 24, 8, 8, 24, 23, 18, 11, 20, 15, 14, 15, 18, 13, 23, 22, 10, 9, 24, 24, 10, 9, 13, 6, 23, 13, 13, 10, 10, 9, 8, 22, 8, 8, 9, 24, 24, 22, 15, 14, 15, 13, 6, 21, 20, 8, 21, 20, 19, 13, 23, 11, 9, 6, 18, 23, 21, 9, 19, 11, 6, 24, 23, 20, 23, 20, 15, 17, 21, 8, 11, 13, 19, 16, 23, 9, 4, 11, 13, 19, 6, 6, 9, 8, 14, 17, 6, 20, 11, 13, 23, 6, 15, 15, 13, 6, 9, 9, 9, 6, 13, 9, 23, 18, 23, 8, 17, 17, 23, 24, 15, 24, 9, 20, 6, 19, 8, 8, 9, 8, 9, 13, 19, 21, 19, 15, 6, 15, 9, 9, 23, 22, 16, 9, 10, 8, 24, 8, 19, 9, 6, 18, 8, 9, 20, 21, 14, 15, 17, 13, 19, 21, 20, 21, 4, 6, 24, 22, 24, 10, 10, 13, 19, 4, 23, 14, 9, 22, 24, 10, 4, 8, 21, 15, 9, 8, 8, 8, 8, 11, 9, 23, 20, 19, 11, 9, 13, 14, 13, 11, 11, 8, 9, 11, 20, 11, 15, 21, 6, 22, 23, 9, 15, 15, 6, 15, 14, 18, 9, 9, 21, 9, 10, 13, 17, 13, 21, 19, 13, 21, 21, 24, 8, 17, 8, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 2, 0, 3, 8, 24, 11, 6, 4, 10, 10, 9, 20, 15, 11, 23, 19, 23, 19, 23, 21, 18, 23, 15, 20, 15, 11, 6, 20, 19, 4, 19, 14, 9, 24, 11, 19, 24, 19, 13, 19, 15, 15, 13, 15, 16, 13, 11, 9, 16, 13, 4, 11, 21, 23, 6, 6, 21, 6, 6, 15, 23, 23, 23, 13, 18, 9, 8, 8, 8, 4, 21, 9, 9, 11, 6, 21, 15, 15, 11, 24, 9, 8, 9, 11, 11, 23, 20, 9, 8, 8, 18, 19, 6, 20, 11, 15, 20, 15, 21, 21, 20, 23, 9, 20, 6, 23, 9, 6, 21, 23, 21, 15, 11, 5, 8, 9, 14, 8, 8, 8, 9, 13, 8, 23, 24, 8, 19, 15, 19, 22, 24, 22, 22, 11, 13, 6, 6, 4, 9, 13, 4, 8, 4, 13, 15, 23, 23, 13, 13, 20, 21, 18, 23, 24, 9, 4, 8, 19, 14, 19, 9, 9, 4, 8, 24, 8, 16, 6, 11, 11, 19, 19, 6, 24, 11, 24, 10, 17, 15, 23, 23, 24, 24, 24, 9, 11, 6, 4, 9, 21, 13, 19, 6, 22, 9, 11, 20, 9, 9, 9, 23, 15, 19, 20, 16, 22, 6, 11, 13, 17, 14, 15, 15, 13, 13, 9, 21, 22, 4, 11, 17, 19, 21, 15, 11, 14, 15, 23, 8, 5, 4, 0, 2, 2, 2, 2),
		(2, 2, 2, 2, 1, 0, 3, 8, 24, 15, 6, 9, 5, 11, 15, 17, 19, 18, 21, 19, 18, 14, 21, 19, 17, 15, 15, 11, 15, 19, 17, 6, 19, 14, 14, 9, 10, 4, 24, 13, 4, 4, 4, 19, 17, 13, 11, 17, 10, 8, 9, 8, 23, 3, 9, 18, 23, 11, 8, 23, 23, 8, 21, 6, 8, 8, 15, 14, 16, 24, 4, 4, 8, 9, 6, 6, 6, 17, 23, 23, 14, 15, 11, 24, 8, 10, 23, 23, 9, 8, 20, 23, 24, 24, 22, 11, 21, 9, 19, 18, 15, 6, 11, 19, 21, 11, 20, 23, 20, 21, 9, 20, 23, 6, 6, 14, 20, 8, 8, 29, 27, 28, 23, 8, 8, 6, 21, 20, 23, 22, 22, 6, 11, 8, 10, 8, 22, 13, 6, 19, 11, 8, 4, 8, 24, 24, 6, 17, 13, 15, 11, 6, 23, 19, 21, 4, 24, 22, 8, 10, 9, 23, 6, 19, 14, 19, 24, 8, 8, 24, 24, 10, 13, 13, 6, 21, 6, 6, 6, 15, 19, 15, 20, 8, 9, 24, 9, 8, 10, 4, 9, 6, 13, 13, 4, 4, 20, 22, 24, 22, 24, 9, 11, 23, 11, 20, 6, 9, 23, 24, 9, 15, 14, 14, 14, 17, 11, 4, 23, 15, 23, 22, 22, 19, 11, 14, 19, 13, 15, 15, 14, 11, 24, 17, 10, 0, 1, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 18, 14, 15, 14, 17, 20, 15, 6, 23, 11, 19, 15, 19, 13, 11, 15, 9, 23, 8, 9, 19, 21, 4, 10, 10, 8, 19, 4, 9, 24, 8, 6, 24, 6, 13, 6, 17, 14, 21, 23, 11, 4, 6, 19, 20, 6, 10, 22, 9, 8, 24, 22, 6, 6, 19, 8, 10, 4, 11, 14, 9, 11, 24, 4, 4, 6, 13, 6, 15, 19, 11, 9, 6, 15, 11, 8, 9, 8, 20, 19, 9, 6, 20, 23, 4, 9, 20, 13, 9, 6, 14, 15, 6, 13, 9, 23, 13, 14, 21, 20, 11, 11, 20, 20, 11, 8, 11, 19, 9, 24, 4, 16, 25, 26, 27, 15, 15, 6, 17, 21, 8, 8, 6, 4, 19, 8, 10, 8, 8, 9, 13, 4, 20, 15, 6, 23, 18, 6, 13, 18, 23, 9, 6, 4, 8, 22, 22, 16, 6, 20, 23, 8, 8, 20, 4, 9, 4, 13, 15, 18, 19, 15, 23, 4, 9, 13, 15, 21, 21, 21, 13, 11, 11, 20, 20, 8, 9, 8, 10, 8, 8, 24, 22, 19, 4, 9, 8, 4, 9, 9, 18, 13, 21, 20, 11, 20, 21, 13, 24, 4, 13, 13, 6, 13, 15, 14, 18, 13, 17, 15, 17, 17, 14, 15, 19, 19, 11, 11, 19, 19, 15, 21, 22, 21, 17, 17, 11, 10, 0, 1, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 18, 13, 6, 11, 11, 11, 11, 21, 15, 15, 21, 13, 4, 9, 23, 9, 11, 23, 8, 4, 11, 15, 9, 13, 9, 4, 6, 8, 10, 4, 3, 9, 22, 13, 13, 17, 14, 13, 23, 13, 9, 8, 20, 14, 13, 6, 8, 8, 10, 10, 10, 9, 9, 19, 18, 9, 8, 6, 21, 11, 8, 4, 9, 4, 6, 19, 6, 13, 13, 6, 20, 9, 11, 15, 11, 6, 6, 6, 14, 13, 6, 23, 8, 23, 11, 10, 9, 19, 19, 4, 19, 14, 10, 11, 20, 21, 18, 21, 19, 23, 20, 18, 11, 13, 6, 6, 23, 11, 6, 10, 8, 16, 25, 26, 27, 15, 18, 19, 6, 6, 8, 23, 6, 20, 21, 4, 8, 10, 10, 9, 15, 23, 23, 21, 20, 8, 20, 4, 9, 15, 15, 23, 6, 8, 8, 8, 10, 8, 11, 19, 23, 9, 20, 23, 24, 11, 9, 16, 13, 15, 14, 19, 23, 11, 18, 9, 9, 11, 11, 21, 19, 11, 4, 23, 20, 23, 8, 8, 8, 8, 24, 22, 6, 24, 4, 6, 6, 8, 6, 11, 11, 11, 14, 15, 21, 18, 15, 13, 24, 11, 17, 17, 14, 14, 15, 13, 23, 11, 6, 17, 13, 11, 11, 11, 14, 19, 13, 13, 6, 14, 13, 4, 8, 11, 15, 15, 13, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 10, 4, 6, 4, 9, 13, 6, 11, 15, 19, 24, 8, 9, 9, 9, 4, 6, 11, 23, 9, 8, 13, 6, 24, 11, 15, 15, 4, 9, 3, 8, 9, 11, 4, 4, 6, 19, 13, 19, 15, 15, 13, 9, 15, 15, 11, 10, 22, 10, 10, 10, 8, 4, 19, 11, 9, 6, 20, 20, 20, 13, 13, 9, 22, 19, 9, 10, 10, 8, 10, 4, 13, 13, 13, 14, 6, 19, 20, 6, 6, 4, 21, 19, 21, 6, 4, 10, 6, 4, 20, 13, 21, 19, 23, 23, 15, 19, 13, 20, 13, 20, 23, 15, 11, 6, 23, 13, 23, 9, 4, 9, 11, 15, 29, 26, 27, 11, 20, 8, 8, 20, 6, 13, 11, 13, 13, 11, 23, 24, 22, 20, 11, 13, 9, 8, 11, 6, 6, 11, 15, 20, 8, 23, 22, 9, 8, 10, 8, 9, 11, 13, 21, 11, 13, 23, 16, 19, 19, 9, 13, 19, 9, 8, 11, 21, 9, 4, 6, 14, 11, 9, 11, 21, 18, 4, 6, 15, 11, 9, 9, 8, 8, 8, 4, 9, 9, 6, 6, 23, 11, 21, 13, 21, 14, 14, 15, 18, 19, 23, 8, 23, 13, 14, 14, 19, 6, 8, 9, 8, 9, 19, 11, 9, 11, 6, 19, 14, 19, 11, 19, 20, 13, 9, 9, 6, 15, 14, 15, 3, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 3, 8, 24, 22, 16, 22, 21, 14, 21, 9, 8, 8, 8, 8, 10, 8, 15, 22, 24, 24, 22, 19, 24, 22, 9, 22, 24, 22, 16, 15, 24, 9, 22, 8, 23, 23, 9, 8, 23, 8, 9, 21, 14, 15, 20, 20, 22, 16, 8, 8, 24, 24, 22, 22, 9, 9, 21, 16, 23, 15, 19, 23, 22, 22, 24, 10, 8, 8, 8, 8, 10, 23, 22, 19, 16, 9, 22, 24, 15, 22, 24, 21, 24, 22, 24, 21, 8, 22, 10, 23, 21, 15, 23, 18, 18, 16, 9, 11, 6, 24, 22, 15, 22, 21, 24, 21, 20, 23, 21, 23, 18, 14, 17, 16, 20, 20, 22, 8, 3, 8, 9, 17, 19, 19, 21, 21, 9, 24, 24, 9, 24, 23, 13, 19, 9, 8, 22, 18, 14, 13, 9, 8, 24, 15, 22, 8, 24, 8, 24, 19, 23, 11, 15, 11, 4, 8, 8, 8, 24, 15, 20, 20, 20, 15, 19, 16, 9, 4, 21, 21, 18, 23, 18, 15, 16, 15, 19, 15, 6, 8, 8, 8, 24, 24, 8, 22, 22, 24, 9, 9, 21, 21, 21, 13, 21, 16, 19, 20, 9, 24, 22, 21, 14, 16, 8, 8, 8, 8, 9, 23, 22, 8, 16, 22, 22, 19, 14, 13, 15, 9, 24, 18, 15, 15, 19, 19, 14, 19, 10, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 0, 12, 4, 22, 22, 24, 22, 17, 17, 23, 8, 4, 10, 8, 22, 9, 11, 8, 8, 8, 6, 19, 17, 13, 11, 19, 20, 9, 11, 13, 15, 11, 11, 14, 13, 22, 24, 10, 8, 24, 3, 9, 11, 19, 14, 6, 20, 17, 13, 17, 17, 13, 22, 11, 6, 11, 13, 19, 11, 13, 15, 4, 10, 9, 11, 6, 10, 8, 23, 8, 8, 6, 9, 11, 17, 11, 9, 9, 6, 17, 9, 13, 6, 13, 13, 6, 11, 11, 19, 17, 17, 9, 17, 17, 15, 11, 16, 11, 24, 11, 13, 6, 14, 6, 6, 17, 17, 17, 17, 13, 17, 19, 13, 9, 22, 19, 15, 5, 8, 8, 4, 11, 15, 11, 22, 15, 24, 10, 9, 8, 9, 21, 24, 9, 16, 6, 11, 13, 14, 17, 17, 13, 11, 6, 6, 17, 13, 8, 10, 24, 24, 6, 11, 9, 13, 13, 17, 13, 13, 14, 11, 6, 11, 13, 17, 17, 17, 15, 23, 21, 18, 19, 6, 15, 15, 18, 15, 13, 11, 17, 8, 10, 8, 10, 8, 10, 9, 9, 10, 8, 24, 13, 23, 9, 19, 6, 11, 6, 11, 13, 17, 13, 15, 17, 8, 8, 8, 8, 6, 11, 11, 19, 11, 11, 9, 9, 15, 14, 14, 17, 17, 5, 23, 5, 11, 11, 14, 14, 19, 12, 0, 0, 1, 1, 1),
		(0, 1, 1, 1, 1, 1, 0, 12, 10, 10, 4, 4, 25, 29, 3, 3, 3, 3, 3, 10, 8, 3, 3, 3, 3, 10, 10, 4, 3, 3, 10, 10, 3, 3, 3, 3, 8, 4, 4, 3, 8, 10, 3, 10, 3, 3, 3, 3, 3, 3, 10, 6, 3, 3, 8, 4, 10, 4, 10, 4, 9, 4, 3, 3, 10, 10, 3, 3, 3, 3, 3, 3, 10, 10, 3, 3, 3, 3, 4, 4, 3, 3, 3, 10, 3, 3, 10, 10, 3, 3, 3, 3, 10, 9, 4, 3, 3, 10, 3, 4, 4, 10, 4, 3, 3, 10, 10, 8, 10, 10, 4, 4, 8, 3, 10, 3, 3, 3, 3, 4, 4, 10, 5, 3, 3, 3, 8, 10, 3, 3, 8, 3, 3, 3, 3, 3, 10, 10, 10, 10, 4, 10, 9, 4, 4, 5, 4, 3, 3, 3, 3, 3, 3, 3, 3, 3, 10, 3, 3, 3, 10, 8, 10, 10, 10, 10, 10, 10, 10, 10, 10, 3, 10, 4, 6, 6, 8, 4, 3, 3, 3, 10, 10, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 10, 3, 3, 10, 3, 3, 4, 6, 10, 3, 3, 3, 3, 3, 10, 10, 10, 10, 3, 3, 3, 4, 4, 4, 4, 3, 3, 10, 29, 3, 10, 4, 4, 4, 3, 0, 1, 1, 1, 1, 1),
		(0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1),
		(0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1),
		(0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1),
		(0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1),
		(0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1),
		(0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1)
	);

	
	signal cor_indice : integer := 0;
	type cor_int is array(0 to 2) of integer range 0 to 255;
	type matriz_cores is array(0 to N_CORES-1) of cor_int;
	constant table_cores: matriz_cores :=
	(
		(164, 167, 170),
		(78, 78, 81),
		(171, 103, 48),
		(219, 224, 232),
		(227, 232, 238),
		(228, 238, 241),
		(233, 237, 243),
		(240, 236, 239),
		(227, 233, 242),
		(231, 235, 243),
		(223, 230, 237),
		(235, 239, 245),
		(214, 210, 216),
		(237, 241, 247),
		(244, 248, 253),
		(241, 245, 251),
		(234, 244, 250),
		(239, 243, 247),
		(239, 243, 251),
		(239, 243, 249),
		(235, 239, 247),
		(237, 241, 249),
		(233, 240, 247),
		(233, 237, 245),
		(230, 237, 245),
		(230, 214, 218),
		(199, 118, 122),
		(212, 162, 166),
		(222, 194, 197),
		(235, 226, 230)
	);



	
	signal pix_x: unsigned(9 downto 0) := unsigned( pixel_x );
	signal pix_y: unsigned(9 downto 0) := unsigned( pixel_y );
	
	begin
	
		pix_x <= unsigned( pixel_x );
		pix_y <= unsigned( pixel_y );

		process( pix_x, pix_y, cor_indice )
		begin
			table_on		 <= '0';
			table_RGB(0) <= "00000000";
			table_RGB(1) <= "00000000";
			table_RGB(2) <= "00000000";
			cor_indice	 <= 0;
			
			if( (Table_Xmin <= pix_x) and (pix_x <= Table_Xmax) and
				 (Table_Ymin <= pix_y) and (pix_y <= Table_Ymax) ) then
				 table_on <= '1';
				 
				 cor_indice   <= table_matriz( img_row_index(  pix_y , Table_Ymin , Table_Ymax, LINHAS ) )
													  ( img_color_index(pix_x , Table_Xmin , Table_Xmax, COLUNAS) );
													  
				 table_RGB(0) <= RGB_UNSIGNED( table_cores(cor_indice)(0) );
				 table_RGB(1) <= RGB_UNSIGNED( table_cores(cor_indice)(1) );
				 table_RGB(2) <= RGB_UNSIGNED( table_cores(cor_indice)(2) );
				 
			end if;
			
		end process;
		
end arch;